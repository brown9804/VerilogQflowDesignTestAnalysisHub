// -----------------------------------------------
// Sumador completo de un bit
// -----------------------------------------------
// Entradas: A, B, Cin
// Salida Cout y S


module sumador_completo (a, b, ci, s, co);
  parameter
    PwrC = 0;

endmodule


// -----------------------------------------------
// Sumador rizado de 8 bits
// -----------------------------------------------
module SUM_RIZADO(a, b, ci, s, co);
  parameter
    PwrC = 0;


endmodule
