module counter_b32 (b32_enable, b32_clk, b32_reset, b32_mode, b32_D, b32_load, b32_rco, b32_Q);

input b32_enable;
input b32_clk;
input b32_reset;
input [1:0] b32_mode;
input [31:0] b32_D;
output [7:0] b32_load;
output [7:0] b32_rco;
output [31:0] b32_Q;

wire vdd = 1'b1;
wire gnd = 1'b0;

	BUFX4 BUFX4_1 ( .A(b32_mode[0]), .Y(b32_mode_0_bF_buf4) );
	BUFX4 BUFX4_2 ( .A(b32_mode[0]), .Y(b32_mode_0_bF_buf3) );
	BUFX4 BUFX4_3 ( .A(b32_mode[0]), .Y(b32_mode_0_bF_buf2) );
	BUFX4 BUFX4_4 ( .A(b32_mode[0]), .Y(b32_mode_0_bF_buf1) );
	BUFX4 BUFX4_5 ( .A(b32_mode[0]), .Y(b32_mode_0_bF_buf0) );
	BUFX4 BUFX4_6 ( .A(b32_clk), .Y(b32_clk_bF_buf7) );
	BUFX4 BUFX4_7 ( .A(b32_clk), .Y(b32_clk_bF_buf6) );
	BUFX4 BUFX4_8 ( .A(b32_clk), .Y(b32_clk_bF_buf5) );
	BUFX4 BUFX4_9 ( .A(b32_clk), .Y(b32_clk_bF_buf4) );
	BUFX4 BUFX4_10 ( .A(b32_clk), .Y(b32_clk_bF_buf3) );
	BUFX4 BUFX4_11 ( .A(b32_clk), .Y(b32_clk_bF_buf2) );
	BUFX4 BUFX4_12 ( .A(b32_clk), .Y(b32_clk_bF_buf1) );
	BUFX4 BUFX4_13 ( .A(b32_clk), .Y(b32_clk_bF_buf0) );
	BUFX4 BUFX4_14 ( .A(b32_mode[1]), .Y(b32_mode_1_bF_buf4) );
	BUFX4 BUFX4_15 ( .A(b32_mode[1]), .Y(b32_mode_1_bF_buf3) );
	BUFX4 BUFX4_16 ( .A(b32_mode[1]), .Y(b32_mode_1_bF_buf2) );
	BUFX4 BUFX4_17 ( .A(b32_mode[1]), .Y(b32_mode_1_bF_buf1) );
	BUFX4 BUFX4_18 ( .A(b32_mode[1]), .Y(b32_mode_1_bF_buf0) );
	DFFPOSX1 DFFPOSX1_1 ( .CLK(b32_clk_bF_buf7), .D(_340__3_), .Q(_0__7_) );
	INVX1 INVX1_1 ( .A(b32_enable), .Y(_397_) );
	NOR2X1 NOR2X1_1 ( .A(b32_reset), .B(_397_), .Y(_398_) );
	INVX4 INVX4_1 ( .A(_398_), .Y(_399_) );
	OAI21X1 OAI21X1_1 ( .A(b32_reset), .B(_397_), .C(_0__8_), .Y(_400_) );
	NAND2X1 NAND2X1_1 ( .A(b32_mode_0_bF_buf4), .B(b32_mode_1_bF_buf4), .Y(_401_) );
	INVX1 INVX1_2 ( .A(b32_mode_0_bF_buf3), .Y(_402_) );
	INVX1 INVX1_3 ( .A(b32_mode_1_bF_buf3), .Y(_403_) );
	OAI21X1 OAI21X1_2 ( .A(_402_), .B(_403_), .C(_0__8_), .Y(_404_) );
	OAI21X1 OAI21X1_3 ( .A(b32_D[8]), .B(_401_), .C(_404_), .Y(_405_) );
	OAI21X1 OAI21X1_4 ( .A(_399_), .B(_405_), .C(_400_), .Y(_396__0_) );
	INVX1 INVX1_4 ( .A(_0__9_), .Y(_406_) );
	INVX1 INVX1_5 ( .A(_401_), .Y(_407_) );
	NOR2X1 NOR2X1_2 ( .A(_0__8_), .B(_0__9_), .Y(_408_) );
	INVX1 INVX1_6 ( .A(_0__8_), .Y(_409_) );
	NOR2X1 NOR2X1_3 ( .A(_409_), .B(_406_), .Y(_410_) );
	OR2X2 OR2X2_1 ( .A(_410_), .B(_408_), .Y(_411_) );
	NOR2X1 NOR2X1_4 ( .A(b32_mode_1_bF_buf2), .B(_402_), .Y(_412_) );
	AOI22X1 AOI22X1_1 ( .A(b32_D[9]), .B(_407_), .C(_412_), .D(_411_), .Y(_413_) );
	NOR2X1 NOR2X1_5 ( .A(_408_), .B(_410_), .Y(_414_) );
	AOI21X1 AOI21X1_1 ( .A(_414_), .B(_402_), .C(_399_), .Y(_415_) );
	AOI22X1 AOI22X1_2 ( .A(_406_), .B(_399_), .C(_415_), .D(_413_), .Y(_396__1_) );
	INVX2 INVX2_1 ( .A(_0__10_), .Y(_416_) );
	NOR2X1 NOR2X1_6 ( .A(b32_mode_0_bF_buf2), .B(_403_), .Y(_417_) );
	NAND3X1 NAND3X1_1 ( .A(_0__8_), .B(_0__9_), .C(_0__10_), .Y(_418_) );
	INVX1 INVX1_7 ( .A(_418_), .Y(_419_) );
	AOI21X1 AOI21X1_2 ( .A(_0__8_), .B(_0__9_), .C(_0__10_), .Y(_420_) );
	OR2X2 OR2X2_2 ( .A(_419_), .B(_420_), .Y(_421_) );
	INVX1 INVX1_8 ( .A(b32_D[10]), .Y(_422_) );
	OAI21X1 OAI21X1_5 ( .A(_422_), .B(_401_), .C(_398_), .Y(_423_) );
	AOI21X1 AOI21X1_3 ( .A(_421_), .B(_417_), .C(_423_), .Y(_424_) );
	NOR2X1 NOR2X1_7 ( .A(b32_mode_0_bF_buf1), .B(b32_mode_1_bF_buf1), .Y(_425_) );
	NOR2X1 NOR2X1_8 ( .A(_420_), .B(_419_), .Y(_426_) );
	NAND2X1 NAND2X1_2 ( .A(_416_), .B(_408_), .Y(_427_) );
	OAI21X1 OAI21X1_6 ( .A(_0__8_), .B(_0__9_), .C(_0__10_), .Y(_428_) );
	NAND2X1 NAND2X1_3 ( .A(_428_), .B(_427_), .Y(_429_) );
	AOI22X1 AOI22X1_3 ( .A(_429_), .B(_412_), .C(_425_), .D(_426_), .Y(_430_) );
	AOI22X1 AOI22X1_4 ( .A(_416_), .B(_399_), .C(_430_), .D(_424_), .Y(_396__2_) );
	INVX4 INVX4_2 ( .A(_0__11_), .Y(_431_) );
	NOR2X1 NOR2X1_9 ( .A(_431_), .B(_418_), .Y(_432_) );
	INVX1 INVX1_9 ( .A(_432_), .Y(_433_) );
	INVX1 INVX1_10 ( .A(_425_), .Y(_434_) );
	AOI21X1 AOI21X1_4 ( .A(_431_), .B(_418_), .C(_434_), .Y(_435_) );
	INVX1 INVX1_11 ( .A(b32_D[11]), .Y(_436_) );
	OAI21X1 OAI21X1_7 ( .A(_436_), .B(_401_), .C(_398_), .Y(_437_) );
	AOI21X1 AOI21X1_5 ( .A(_433_), .B(_435_), .C(_437_), .Y(_438_) );
	NAND3X1 NAND3X1_2 ( .A(_416_), .B(_431_), .C(_408_), .Y(_439_) );
	OR2X2 OR2X2_3 ( .A(_0__8_), .B(_0__9_), .Y(_440_) );
	OAI21X1 OAI21X1_8 ( .A(_0__10_), .B(_440_), .C(_0__11_), .Y(_441_) );
	NAND2X1 NAND2X1_4 ( .A(_439_), .B(_441_), .Y(_442_) );
	XNOR2X1 XNOR2X1_1 ( .A(_420_), .B(_431_), .Y(_443_) );
	AOI22X1 AOI22X1_5 ( .A(_417_), .B(_443_), .C(_412_), .D(_442_), .Y(_444_) );
	AOI22X1 AOI22X1_6 ( .A(_431_), .B(_399_), .C(_438_), .D(_444_), .Y(_396__3_) );
	NOR2X1 NOR2X1_10 ( .A(_409_), .B(_399_), .Y(_393__0_) );
	NOR2X1 NOR2X1_11 ( .A(_406_), .B(_399_), .Y(_393__1_) );
	NOR2X1 NOR2X1_12 ( .A(_416_), .B(_399_), .Y(_393__2_) );
	NOR2X1 NOR2X1_13 ( .A(_431_), .B(_399_), .Y(_393__3_) );
	INVX1 INVX1_12 ( .A(_439_), .Y(_445_) );
	NAND2X1 NAND2X1_5 ( .A(_412_), .B(_445_), .Y(_446_) );
	AND2X2 AND2X2_1 ( .A(_420_), .B(_431_), .Y(_447_) );
	AOI22X1 AOI22X1_7 ( .A(_425_), .B(_432_), .C(_417_), .D(_447_), .Y(_448_) );
	AOI21X1 AOI21X1_6 ( .A(_446_), .B(_448_), .C(_399_), .Y(_395_) );
	NOR2X1 NOR2X1_14 ( .A(_401_), .B(_399_), .Y(_394_) );
	DFFPOSX1 DFFPOSX1_2 ( .CLK(b32_clk_bF_buf6), .D(_394_), .Q(counter_8b11_b4_load) );
	DFFPOSX1 DFFPOSX1_3 ( .CLK(b32_clk_bF_buf5), .D(_395_), .Q(counter_8b11_b4_rco) );
	DFFPOSX1 DFFPOSX1_4 ( .CLK(b32_clk_bF_buf4), .D(_393__0_), .Q(_0__8_) );
	DFFPOSX1 DFFPOSX1_5 ( .CLK(b32_clk_bF_buf3), .D(_393__1_), .Q(_0__9_) );
	DFFPOSX1 DFFPOSX1_6 ( .CLK(b32_clk_bF_buf2), .D(_393__2_), .Q(_0__10_) );
	DFFPOSX1 DFFPOSX1_7 ( .CLK(b32_clk_bF_buf1), .D(_393__3_), .Q(_0__11_) );
	DFFPOSX1 DFFPOSX1_8 ( .CLK(b32_clk_bF_buf0), .D(_396__0_), .Q(_0__8_) );
	DFFPOSX1 DFFPOSX1_9 ( .CLK(b32_clk_bF_buf7), .D(_396__1_), .Q(_0__9_) );
	DFFPOSX1 DFFPOSX1_10 ( .CLK(b32_clk_bF_buf6), .D(_396__2_), .Q(_0__10_) );
	DFFPOSX1 DFFPOSX1_11 ( .CLK(b32_clk_bF_buf5), .D(_396__3_), .Q(_0__11_) );
	BUFX2 BUFX2_1 ( .A(_0__0_), .Y(b32_Q[0]) );
	BUFX2 BUFX2_2 ( .A(_0__1_), .Y(b32_Q[1]) );
	BUFX2 BUFX2_3 ( .A(_0__2_), .Y(b32_Q[2]) );
	BUFX2 BUFX2_4 ( .A(_0__3_), .Y(b32_Q[3]) );
	BUFX2 BUFX2_5 ( .A(_0__4_), .Y(b32_Q[4]) );
	BUFX2 BUFX2_6 ( .A(_0__5_), .Y(b32_Q[5]) );
	BUFX2 BUFX2_7 ( .A(_0__6_), .Y(b32_Q[6]) );
	BUFX2 BUFX2_8 ( .A(_0__7_), .Y(b32_Q[7]) );
	BUFX2 BUFX2_9 ( .A(_0__8_), .Y(b32_Q[8]) );
	BUFX2 BUFX2_10 ( .A(_0__9_), .Y(b32_Q[9]) );
	BUFX2 BUFX2_11 ( .A(_0__10_), .Y(b32_Q[10]) );
	BUFX2 BUFX2_12 ( .A(_0__11_), .Y(b32_Q[11]) );
	BUFX2 BUFX2_13 ( .A(_0__12_), .Y(b32_Q[12]) );
	BUFX2 BUFX2_14 ( .A(_0__13_), .Y(b32_Q[13]) );
	BUFX2 BUFX2_15 ( .A(_0__14_), .Y(b32_Q[14]) );
	BUFX2 BUFX2_16 ( .A(_0__15_), .Y(b32_Q[15]) );
	BUFX2 BUFX2_17 ( .A(_0__16_), .Y(b32_Q[16]) );
	BUFX2 BUFX2_18 ( .A(_0__17_), .Y(b32_Q[17]) );
	BUFX2 BUFX2_19 ( .A(_0__18_), .Y(b32_Q[18]) );
	BUFX2 BUFX2_20 ( .A(_0__19_), .Y(b32_Q[19]) );
	BUFX2 BUFX2_21 ( .A(_0__20_), .Y(b32_Q[20]) );
	BUFX2 BUFX2_22 ( .A(_0__21_), .Y(b32_Q[21]) );
	BUFX2 BUFX2_23 ( .A(_0__22_), .Y(b32_Q[22]) );
	BUFX2 BUFX2_24 ( .A(_0__23_), .Y(b32_Q[23]) );
	BUFX2 BUFX2_25 ( .A(_0__24_), .Y(b32_Q[24]) );
	BUFX2 BUFX2_26 ( .A(_0__25_), .Y(b32_Q[25]) );
	BUFX2 BUFX2_27 ( .A(_0__26_), .Y(b32_Q[26]) );
	BUFX2 BUFX2_28 ( .A(_0__27_), .Y(b32_Q[27]) );
	BUFX2 BUFX2_29 ( .A(_0__28_), .Y(b32_Q[28]) );
	BUFX2 BUFX2_30 ( .A(_0__29_), .Y(b32_Q[29]) );
	BUFX2 BUFX2_31 ( .A(_0__30_), .Y(b32_Q[30]) );
	BUFX2 BUFX2_32 ( .A(_0__31_), .Y(b32_Q[31]) );
	BUFX2 BUFX2_33 ( .A(counter_0b3_b4_load), .Y(b32_load[0]) );
	BUFX2 BUFX2_34 ( .A(counter_4b7_b4_load), .Y(b32_load[1]) );
	BUFX2 BUFX2_35 ( .A(counter_8b11_b4_load), .Y(b32_load[2]) );
	BUFX2 BUFX2_36 ( .A(counter_12b15_b4_load), .Y(b32_load[3]) );
	BUFX2 BUFX2_37 ( .A(counter_16b19_b4_load), .Y(b32_load[4]) );
	BUFX2 BUFX2_38 ( .A(counter_20b23_b4_load), .Y(b32_load[5]) );
	BUFX2 BUFX2_39 ( .A(counter_24b27_b4_load), .Y(b32_load[6]) );
	BUFX2 BUFX2_40 ( .A(counter_28b31_b4_load), .Y(b32_load[7]) );
	BUFX2 BUFX2_41 ( .A(counter_0b3_b4_rco), .Y(b32_rco[0]) );
	BUFX2 BUFX2_42 ( .A(counter_4b7_b4_rco), .Y(b32_rco[1]) );
	BUFX2 BUFX2_43 ( .A(counter_8b11_b4_rco), .Y(b32_rco[2]) );
	BUFX2 BUFX2_44 ( .A(counter_12b15_b4_rco), .Y(b32_rco[3]) );
	BUFX2 BUFX2_45 ( .A(counter_16b19_b4_rco), .Y(b32_rco[4]) );
	BUFX2 BUFX2_46 ( .A(counter_20b23_b4_rco), .Y(b32_rco[5]) );
	BUFX2 BUFX2_47 ( .A(counter_24b27_b4_rco), .Y(b32_rco[6]) );
	BUFX2 BUFX2_48 ( .A(counter_28b31_b4_rco), .Y(b32_rco[7]) );
	INVX1 INVX1_13 ( .A(b32_enable), .Y(_5_) );
	NOR2X1 NOR2X1_15 ( .A(b32_reset), .B(_5_), .Y(_6_) );
	INVX4 INVX4_3 ( .A(_6_), .Y(_7_) );
	OAI21X1 OAI21X1_9 ( .A(b32_reset), .B(_5_), .C(_0__0_), .Y(_8_) );
	NAND2X1 NAND2X1_6 ( .A(b32_mode_0_bF_buf0), .B(b32_mode_1_bF_buf0), .Y(_9_) );
	INVX1 INVX1_14 ( .A(b32_mode_0_bF_buf4), .Y(_10_) );
	INVX1 INVX1_15 ( .A(b32_mode_1_bF_buf4), .Y(_11_) );
	OAI21X1 OAI21X1_10 ( .A(_10_), .B(_11_), .C(_0__0_), .Y(_12_) );
	OAI21X1 OAI21X1_11 ( .A(b32_D[0]), .B(_9_), .C(_12_), .Y(_13_) );
	OAI21X1 OAI21X1_12 ( .A(_7_), .B(_13_), .C(_8_), .Y(_4__0_) );
	INVX1 INVX1_16 ( .A(_0__1_), .Y(_14_) );
	INVX1 INVX1_17 ( .A(_9_), .Y(_15_) );
	NOR2X1 NOR2X1_16 ( .A(_0__0_), .B(_0__1_), .Y(_16_) );
	INVX1 INVX1_18 ( .A(_0__0_), .Y(_17_) );
	NOR2X1 NOR2X1_17 ( .A(_17_), .B(_14_), .Y(_18_) );
	OR2X2 OR2X2_4 ( .A(_18_), .B(_16_), .Y(_19_) );
	NOR2X1 NOR2X1_18 ( .A(b32_mode_1_bF_buf3), .B(_10_), .Y(_20_) );
	AOI22X1 AOI22X1_8 ( .A(b32_D[1]), .B(_15_), .C(_20_), .D(_19_), .Y(_21_) );
	NOR2X1 NOR2X1_19 ( .A(_16_), .B(_18_), .Y(_22_) );
	AOI21X1 AOI21X1_7 ( .A(_22_), .B(_10_), .C(_7_), .Y(_23_) );
	AOI22X1 AOI22X1_9 ( .A(_14_), .B(_7_), .C(_23_), .D(_21_), .Y(_4__1_) );
	INVX2 INVX2_2 ( .A(_0__2_), .Y(_24_) );
	NOR2X1 NOR2X1_20 ( .A(b32_mode_0_bF_buf3), .B(_11_), .Y(_25_) );
	NAND3X1 NAND3X1_3 ( .A(_0__0_), .B(_0__1_), .C(_0__2_), .Y(_26_) );
	INVX1 INVX1_19 ( .A(_26_), .Y(_27_) );
	AOI21X1 AOI21X1_8 ( .A(_0__0_), .B(_0__1_), .C(_0__2_), .Y(_28_) );
	OR2X2 OR2X2_5 ( .A(_27_), .B(_28_), .Y(_29_) );
	INVX1 INVX1_20 ( .A(b32_D[2]), .Y(_30_) );
	OAI21X1 OAI21X1_13 ( .A(_30_), .B(_9_), .C(_6_), .Y(_31_) );
	AOI21X1 AOI21X1_9 ( .A(_29_), .B(_25_), .C(_31_), .Y(_32_) );
	NOR2X1 NOR2X1_21 ( .A(b32_mode_0_bF_buf2), .B(b32_mode_1_bF_buf2), .Y(_33_) );
	NOR2X1 NOR2X1_22 ( .A(_28_), .B(_27_), .Y(_34_) );
	NAND2X1 NAND2X1_7 ( .A(_24_), .B(_16_), .Y(_35_) );
	OAI21X1 OAI21X1_14 ( .A(_0__0_), .B(_0__1_), .C(_0__2_), .Y(_36_) );
	NAND2X1 NAND2X1_8 ( .A(_36_), .B(_35_), .Y(_37_) );
	AOI22X1 AOI22X1_10 ( .A(_37_), .B(_20_), .C(_33_), .D(_34_), .Y(_38_) );
	AOI22X1 AOI22X1_11 ( .A(_24_), .B(_7_), .C(_38_), .D(_32_), .Y(_4__2_) );
	INVX4 INVX4_4 ( .A(_0__3_), .Y(_39_) );
	NOR2X1 NOR2X1_23 ( .A(_39_), .B(_26_), .Y(_40_) );
	INVX1 INVX1_21 ( .A(_40_), .Y(_41_) );
	INVX1 INVX1_22 ( .A(_33_), .Y(_42_) );
	AOI21X1 AOI21X1_10 ( .A(_39_), .B(_26_), .C(_42_), .Y(_43_) );
	INVX1 INVX1_23 ( .A(b32_D[3]), .Y(_44_) );
	OAI21X1 OAI21X1_15 ( .A(_44_), .B(_9_), .C(_6_), .Y(_45_) );
	AOI21X1 AOI21X1_11 ( .A(_41_), .B(_43_), .C(_45_), .Y(_46_) );
	NAND3X1 NAND3X1_4 ( .A(_24_), .B(_39_), .C(_16_), .Y(_47_) );
	OR2X2 OR2X2_6 ( .A(_0__0_), .B(_0__1_), .Y(_48_) );
	OAI21X1 OAI21X1_16 ( .A(_0__2_), .B(_48_), .C(_0__3_), .Y(_49_) );
	NAND2X1 NAND2X1_9 ( .A(_47_), .B(_49_), .Y(_50_) );
	XNOR2X1 XNOR2X1_2 ( .A(_28_), .B(_39_), .Y(_51_) );
	AOI22X1 AOI22X1_12 ( .A(_25_), .B(_51_), .C(_20_), .D(_50_), .Y(_52_) );
	AOI22X1 AOI22X1_13 ( .A(_39_), .B(_7_), .C(_46_), .D(_52_), .Y(_4__3_) );
	NOR2X1 NOR2X1_24 ( .A(_17_), .B(_7_), .Y(_1__0_) );
	NOR2X1 NOR2X1_25 ( .A(_14_), .B(_7_), .Y(_1__1_) );
	NOR2X1 NOR2X1_26 ( .A(_24_), .B(_7_), .Y(_1__2_) );
	NOR2X1 NOR2X1_27 ( .A(_39_), .B(_7_), .Y(_1__3_) );
	INVX1 INVX1_24 ( .A(_47_), .Y(_53_) );
	NAND2X1 NAND2X1_10 ( .A(_20_), .B(_53_), .Y(_54_) );
	AND2X2 AND2X2_2 ( .A(_28_), .B(_39_), .Y(_55_) );
	AOI22X1 AOI22X1_14 ( .A(_33_), .B(_40_), .C(_25_), .D(_55_), .Y(_56_) );
	AOI21X1 AOI21X1_12 ( .A(_54_), .B(_56_), .C(_7_), .Y(_3_) );
	NOR2X1 NOR2X1_28 ( .A(_9_), .B(_7_), .Y(_2_) );
	DFFPOSX1 DFFPOSX1_12 ( .CLK(b32_clk_bF_buf4), .D(_2_), .Q(counter_0b3_b4_load) );
	DFFPOSX1 DFFPOSX1_13 ( .CLK(b32_clk_bF_buf3), .D(_3_), .Q(counter_0b3_b4_rco) );
	DFFPOSX1 DFFPOSX1_14 ( .CLK(b32_clk_bF_buf2), .D(_1__0_), .Q(_0__0_) );
	DFFPOSX1 DFFPOSX1_15 ( .CLK(b32_clk_bF_buf1), .D(_1__1_), .Q(_0__1_) );
	DFFPOSX1 DFFPOSX1_16 ( .CLK(b32_clk_bF_buf0), .D(_1__2_), .Q(_0__2_) );
	DFFPOSX1 DFFPOSX1_17 ( .CLK(b32_clk_bF_buf7), .D(_1__3_), .Q(_0__3_) );
	DFFPOSX1 DFFPOSX1_18 ( .CLK(b32_clk_bF_buf6), .D(_4__0_), .Q(_0__0_) );
	DFFPOSX1 DFFPOSX1_19 ( .CLK(b32_clk_bF_buf5), .D(_4__1_), .Q(_0__1_) );
	DFFPOSX1 DFFPOSX1_20 ( .CLK(b32_clk_bF_buf4), .D(_4__2_), .Q(_0__2_) );
	DFFPOSX1 DFFPOSX1_21 ( .CLK(b32_clk_bF_buf3), .D(_4__3_), .Q(_0__3_) );
	INVX1 INVX1_25 ( .A(b32_enable), .Y(_61_) );
	NOR2X1 NOR2X1_29 ( .A(b32_reset), .B(_61_), .Y(_62_) );
	INVX4 INVX4_5 ( .A(_62_), .Y(_63_) );
	OAI21X1 OAI21X1_17 ( .A(b32_reset), .B(_61_), .C(_0__12_), .Y(_64_) );
	NAND2X1 NAND2X1_11 ( .A(b32_mode_0_bF_buf1), .B(b32_mode_1_bF_buf1), .Y(_65_) );
	INVX1 INVX1_26 ( .A(b32_mode_0_bF_buf0), .Y(_66_) );
	INVX1 INVX1_27 ( .A(b32_mode_1_bF_buf0), .Y(_67_) );
	OAI21X1 OAI21X1_18 ( .A(_66_), .B(_67_), .C(_0__12_), .Y(_68_) );
	OAI21X1 OAI21X1_19 ( .A(b32_D[12]), .B(_65_), .C(_68_), .Y(_69_) );
	OAI21X1 OAI21X1_20 ( .A(_63_), .B(_69_), .C(_64_), .Y(_60__0_) );
	INVX1 INVX1_28 ( .A(_0__13_), .Y(_70_) );
	INVX1 INVX1_29 ( .A(_65_), .Y(_71_) );
	NOR2X1 NOR2X1_30 ( .A(_0__12_), .B(_0__13_), .Y(_72_) );
	INVX1 INVX1_30 ( .A(_0__12_), .Y(_73_) );
	NOR2X1 NOR2X1_31 ( .A(_73_), .B(_70_), .Y(_74_) );
	OR2X2 OR2X2_7 ( .A(_74_), .B(_72_), .Y(_75_) );
	NOR2X1 NOR2X1_32 ( .A(b32_mode_1_bF_buf4), .B(_66_), .Y(_76_) );
	AOI22X1 AOI22X1_15 ( .A(b32_D[13]), .B(_71_), .C(_76_), .D(_75_), .Y(_77_) );
	NOR2X1 NOR2X1_33 ( .A(_72_), .B(_74_), .Y(_78_) );
	AOI21X1 AOI21X1_13 ( .A(_78_), .B(_66_), .C(_63_), .Y(_79_) );
	AOI22X1 AOI22X1_16 ( .A(_70_), .B(_63_), .C(_79_), .D(_77_), .Y(_60__1_) );
	INVX2 INVX2_3 ( .A(_0__14_), .Y(_80_) );
	NOR2X1 NOR2X1_34 ( .A(b32_mode_0_bF_buf4), .B(_67_), .Y(_81_) );
	NAND3X1 NAND3X1_5 ( .A(_0__12_), .B(_0__13_), .C(_0__14_), .Y(_82_) );
	INVX1 INVX1_31 ( .A(_82_), .Y(_83_) );
	AOI21X1 AOI21X1_14 ( .A(_0__12_), .B(_0__13_), .C(_0__14_), .Y(_84_) );
	OR2X2 OR2X2_8 ( .A(_83_), .B(_84_), .Y(_85_) );
	INVX1 INVX1_32 ( .A(b32_D[14]), .Y(_86_) );
	OAI21X1 OAI21X1_21 ( .A(_86_), .B(_65_), .C(_62_), .Y(_87_) );
	AOI21X1 AOI21X1_15 ( .A(_85_), .B(_81_), .C(_87_), .Y(_88_) );
	NOR2X1 NOR2X1_35 ( .A(b32_mode_0_bF_buf3), .B(b32_mode_1_bF_buf3), .Y(_89_) );
	NOR2X1 NOR2X1_36 ( .A(_84_), .B(_83_), .Y(_90_) );
	NAND2X1 NAND2X1_12 ( .A(_80_), .B(_72_), .Y(_91_) );
	OAI21X1 OAI21X1_22 ( .A(_0__12_), .B(_0__13_), .C(_0__14_), .Y(_92_) );
	NAND2X1 NAND2X1_13 ( .A(_92_), .B(_91_), .Y(_93_) );
	AOI22X1 AOI22X1_17 ( .A(_93_), .B(_76_), .C(_89_), .D(_90_), .Y(_94_) );
	AOI22X1 AOI22X1_18 ( .A(_80_), .B(_63_), .C(_94_), .D(_88_), .Y(_60__2_) );
	INVX4 INVX4_6 ( .A(_0__15_), .Y(_95_) );
	NOR2X1 NOR2X1_37 ( .A(_95_), .B(_82_), .Y(_96_) );
	INVX1 INVX1_33 ( .A(_96_), .Y(_97_) );
	INVX1 INVX1_34 ( .A(_89_), .Y(_98_) );
	AOI21X1 AOI21X1_16 ( .A(_95_), .B(_82_), .C(_98_), .Y(_99_) );
	INVX1 INVX1_35 ( .A(b32_D[15]), .Y(_100_) );
	OAI21X1 OAI21X1_23 ( .A(_100_), .B(_65_), .C(_62_), .Y(_101_) );
	AOI21X1 AOI21X1_17 ( .A(_97_), .B(_99_), .C(_101_), .Y(_102_) );
	NAND3X1 NAND3X1_6 ( .A(_80_), .B(_95_), .C(_72_), .Y(_103_) );
	OR2X2 OR2X2_9 ( .A(_0__12_), .B(_0__13_), .Y(_104_) );
	OAI21X1 OAI21X1_24 ( .A(_0__14_), .B(_104_), .C(_0__15_), .Y(_105_) );
	NAND2X1 NAND2X1_14 ( .A(_103_), .B(_105_), .Y(_106_) );
	XNOR2X1 XNOR2X1_3 ( .A(_84_), .B(_95_), .Y(_107_) );
	AOI22X1 AOI22X1_19 ( .A(_81_), .B(_107_), .C(_76_), .D(_106_), .Y(_108_) );
	AOI22X1 AOI22X1_20 ( .A(_95_), .B(_63_), .C(_102_), .D(_108_), .Y(_60__3_) );
	NOR2X1 NOR2X1_38 ( .A(_73_), .B(_63_), .Y(_57__0_) );
	NOR2X1 NOR2X1_39 ( .A(_70_), .B(_63_), .Y(_57__1_) );
	NOR2X1 NOR2X1_40 ( .A(_80_), .B(_63_), .Y(_57__2_) );
	NOR2X1 NOR2X1_41 ( .A(_95_), .B(_63_), .Y(_57__3_) );
	INVX1 INVX1_36 ( .A(_103_), .Y(_109_) );
	NAND2X1 NAND2X1_15 ( .A(_76_), .B(_109_), .Y(_110_) );
	AND2X2 AND2X2_3 ( .A(_84_), .B(_95_), .Y(_111_) );
	AOI22X1 AOI22X1_21 ( .A(_89_), .B(_96_), .C(_81_), .D(_111_), .Y(_112_) );
	AOI21X1 AOI21X1_18 ( .A(_110_), .B(_112_), .C(_63_), .Y(_59_) );
	NOR2X1 NOR2X1_42 ( .A(_65_), .B(_63_), .Y(_58_) );
	DFFPOSX1 DFFPOSX1_22 ( .CLK(b32_clk_bF_buf2), .D(_58_), .Q(counter_12b15_b4_load) );
	DFFPOSX1 DFFPOSX1_23 ( .CLK(b32_clk_bF_buf1), .D(_59_), .Q(counter_12b15_b4_rco) );
	DFFPOSX1 DFFPOSX1_24 ( .CLK(b32_clk_bF_buf0), .D(_57__0_), .Q(_0__12_) );
	DFFPOSX1 DFFPOSX1_25 ( .CLK(b32_clk_bF_buf7), .D(_57__1_), .Q(_0__13_) );
	DFFPOSX1 DFFPOSX1_26 ( .CLK(b32_clk_bF_buf6), .D(_57__2_), .Q(_0__14_) );
	DFFPOSX1 DFFPOSX1_27 ( .CLK(b32_clk_bF_buf5), .D(_57__3_), .Q(_0__15_) );
	DFFPOSX1 DFFPOSX1_28 ( .CLK(b32_clk_bF_buf4), .D(_60__0_), .Q(_0__12_) );
	DFFPOSX1 DFFPOSX1_29 ( .CLK(b32_clk_bF_buf3), .D(_60__1_), .Q(_0__13_) );
	DFFPOSX1 DFFPOSX1_30 ( .CLK(b32_clk_bF_buf2), .D(_60__2_), .Q(_0__14_) );
	DFFPOSX1 DFFPOSX1_31 ( .CLK(b32_clk_bF_buf1), .D(_60__3_), .Q(_0__15_) );
	INVX1 INVX1_37 ( .A(b32_enable), .Y(_117_) );
	NOR2X1 NOR2X1_43 ( .A(b32_reset), .B(_117_), .Y(_118_) );
	INVX4 INVX4_7 ( .A(_118_), .Y(_119_) );
	OAI21X1 OAI21X1_25 ( .A(b32_reset), .B(_117_), .C(_0__16_), .Y(_120_) );
	NAND2X1 NAND2X1_16 ( .A(b32_mode_0_bF_buf2), .B(b32_mode_1_bF_buf2), .Y(_121_) );
	INVX1 INVX1_38 ( .A(b32_mode_0_bF_buf1), .Y(_122_) );
	INVX1 INVX1_39 ( .A(b32_mode_1_bF_buf1), .Y(_123_) );
	OAI21X1 OAI21X1_26 ( .A(_122_), .B(_123_), .C(_0__16_), .Y(_124_) );
	OAI21X1 OAI21X1_27 ( .A(b32_D[16]), .B(_121_), .C(_124_), .Y(_125_) );
	OAI21X1 OAI21X1_28 ( .A(_119_), .B(_125_), .C(_120_), .Y(_116__0_) );
	INVX1 INVX1_40 ( .A(_0__17_), .Y(_126_) );
	INVX1 INVX1_41 ( .A(_121_), .Y(_127_) );
	NOR2X1 NOR2X1_44 ( .A(_0__16_), .B(_0__17_), .Y(_128_) );
	INVX1 INVX1_42 ( .A(_0__16_), .Y(_129_) );
	NOR2X1 NOR2X1_45 ( .A(_129_), .B(_126_), .Y(_130_) );
	OR2X2 OR2X2_10 ( .A(_130_), .B(_128_), .Y(_131_) );
	NOR2X1 NOR2X1_46 ( .A(b32_mode_1_bF_buf0), .B(_122_), .Y(_132_) );
	AOI22X1 AOI22X1_22 ( .A(b32_D[17]), .B(_127_), .C(_132_), .D(_131_), .Y(_133_) );
	NOR2X1 NOR2X1_47 ( .A(_128_), .B(_130_), .Y(_134_) );
	AOI21X1 AOI21X1_19 ( .A(_134_), .B(_122_), .C(_119_), .Y(_135_) );
	AOI22X1 AOI22X1_23 ( .A(_126_), .B(_119_), .C(_135_), .D(_133_), .Y(_116__1_) );
	INVX2 INVX2_4 ( .A(_0__18_), .Y(_136_) );
	NOR2X1 NOR2X1_48 ( .A(b32_mode_0_bF_buf0), .B(_123_), .Y(_137_) );
	NAND3X1 NAND3X1_7 ( .A(_0__16_), .B(_0__17_), .C(_0__18_), .Y(_138_) );
	INVX1 INVX1_43 ( .A(_138_), .Y(_139_) );
	AOI21X1 AOI21X1_20 ( .A(_0__16_), .B(_0__17_), .C(_0__18_), .Y(_140_) );
	OR2X2 OR2X2_11 ( .A(_139_), .B(_140_), .Y(_141_) );
	INVX1 INVX1_44 ( .A(b32_D[18]), .Y(_142_) );
	OAI21X1 OAI21X1_29 ( .A(_142_), .B(_121_), .C(_118_), .Y(_143_) );
	AOI21X1 AOI21X1_21 ( .A(_141_), .B(_137_), .C(_143_), .Y(_144_) );
	NOR2X1 NOR2X1_49 ( .A(b32_mode_0_bF_buf4), .B(b32_mode_1_bF_buf4), .Y(_145_) );
	NOR2X1 NOR2X1_50 ( .A(_140_), .B(_139_), .Y(_146_) );
	NAND2X1 NAND2X1_17 ( .A(_136_), .B(_128_), .Y(_147_) );
	OAI21X1 OAI21X1_30 ( .A(_0__16_), .B(_0__17_), .C(_0__18_), .Y(_148_) );
	NAND2X1 NAND2X1_18 ( .A(_148_), .B(_147_), .Y(_149_) );
	AOI22X1 AOI22X1_24 ( .A(_149_), .B(_132_), .C(_145_), .D(_146_), .Y(_150_) );
	AOI22X1 AOI22X1_25 ( .A(_136_), .B(_119_), .C(_150_), .D(_144_), .Y(_116__2_) );
	INVX4 INVX4_8 ( .A(_0__19_), .Y(_151_) );
	NOR2X1 NOR2X1_51 ( .A(_151_), .B(_138_), .Y(_152_) );
	INVX1 INVX1_45 ( .A(_152_), .Y(_153_) );
	INVX1 INVX1_46 ( .A(_145_), .Y(_154_) );
	AOI21X1 AOI21X1_22 ( .A(_151_), .B(_138_), .C(_154_), .Y(_155_) );
	INVX1 INVX1_47 ( .A(b32_D[19]), .Y(_156_) );
	OAI21X1 OAI21X1_31 ( .A(_156_), .B(_121_), .C(_118_), .Y(_157_) );
	AOI21X1 AOI21X1_23 ( .A(_153_), .B(_155_), .C(_157_), .Y(_158_) );
	NAND3X1 NAND3X1_8 ( .A(_136_), .B(_151_), .C(_128_), .Y(_159_) );
	OR2X2 OR2X2_12 ( .A(_0__16_), .B(_0__17_), .Y(_160_) );
	OAI21X1 OAI21X1_32 ( .A(_0__18_), .B(_160_), .C(_0__19_), .Y(_161_) );
	NAND2X1 NAND2X1_19 ( .A(_159_), .B(_161_), .Y(_162_) );
	XNOR2X1 XNOR2X1_4 ( .A(_140_), .B(_151_), .Y(_163_) );
	AOI22X1 AOI22X1_26 ( .A(_137_), .B(_163_), .C(_132_), .D(_162_), .Y(_164_) );
	AOI22X1 AOI22X1_27 ( .A(_151_), .B(_119_), .C(_158_), .D(_164_), .Y(_116__3_) );
	NOR2X1 NOR2X1_52 ( .A(_129_), .B(_119_), .Y(_113__0_) );
	NOR2X1 NOR2X1_53 ( .A(_126_), .B(_119_), .Y(_113__1_) );
	NOR2X1 NOR2X1_54 ( .A(_136_), .B(_119_), .Y(_113__2_) );
	NOR2X1 NOR2X1_55 ( .A(_151_), .B(_119_), .Y(_113__3_) );
	INVX1 INVX1_48 ( .A(_159_), .Y(_165_) );
	NAND2X1 NAND2X1_20 ( .A(_132_), .B(_165_), .Y(_166_) );
	AND2X2 AND2X2_4 ( .A(_140_), .B(_151_), .Y(_167_) );
	AOI22X1 AOI22X1_28 ( .A(_145_), .B(_152_), .C(_137_), .D(_167_), .Y(_168_) );
	AOI21X1 AOI21X1_24 ( .A(_166_), .B(_168_), .C(_119_), .Y(_115_) );
	NOR2X1 NOR2X1_56 ( .A(_121_), .B(_119_), .Y(_114_) );
	DFFPOSX1 DFFPOSX1_32 ( .CLK(b32_clk_bF_buf0), .D(_114_), .Q(counter_16b19_b4_load) );
	DFFPOSX1 DFFPOSX1_33 ( .CLK(b32_clk_bF_buf7), .D(_115_), .Q(counter_16b19_b4_rco) );
	DFFPOSX1 DFFPOSX1_34 ( .CLK(b32_clk_bF_buf6), .D(_113__0_), .Q(_0__16_) );
	DFFPOSX1 DFFPOSX1_35 ( .CLK(b32_clk_bF_buf5), .D(_113__1_), .Q(_0__17_) );
	DFFPOSX1 DFFPOSX1_36 ( .CLK(b32_clk_bF_buf4), .D(_113__2_), .Q(_0__18_) );
	DFFPOSX1 DFFPOSX1_37 ( .CLK(b32_clk_bF_buf3), .D(_113__3_), .Q(_0__19_) );
	DFFPOSX1 DFFPOSX1_38 ( .CLK(b32_clk_bF_buf2), .D(_116__0_), .Q(_0__16_) );
	DFFPOSX1 DFFPOSX1_39 ( .CLK(b32_clk_bF_buf1), .D(_116__1_), .Q(_0__17_) );
	DFFPOSX1 DFFPOSX1_40 ( .CLK(b32_clk_bF_buf0), .D(_116__2_), .Q(_0__18_) );
	DFFPOSX1 DFFPOSX1_41 ( .CLK(b32_clk_bF_buf7), .D(_116__3_), .Q(_0__19_) );
	INVX1 INVX1_49 ( .A(b32_enable), .Y(_173_) );
	NOR2X1 NOR2X1_57 ( .A(b32_reset), .B(_173_), .Y(_174_) );
	INVX4 INVX4_9 ( .A(_174_), .Y(_175_) );
	OAI21X1 OAI21X1_33 ( .A(b32_reset), .B(_173_), .C(_0__20_), .Y(_176_) );
	NAND2X1 NAND2X1_21 ( .A(b32_mode_0_bF_buf3), .B(b32_mode_1_bF_buf3), .Y(_177_) );
	INVX1 INVX1_50 ( .A(b32_mode_0_bF_buf2), .Y(_178_) );
	INVX1 INVX1_51 ( .A(b32_mode_1_bF_buf2), .Y(_179_) );
	OAI21X1 OAI21X1_34 ( .A(_178_), .B(_179_), .C(_0__20_), .Y(_180_) );
	OAI21X1 OAI21X1_35 ( .A(b32_D[20]), .B(_177_), .C(_180_), .Y(_181_) );
	OAI21X1 OAI21X1_36 ( .A(_175_), .B(_181_), .C(_176_), .Y(_172__0_) );
	INVX1 INVX1_52 ( .A(_0__21_), .Y(_182_) );
	INVX1 INVX1_53 ( .A(_177_), .Y(_183_) );
	NOR2X1 NOR2X1_58 ( .A(_0__20_), .B(_0__21_), .Y(_184_) );
	INVX1 INVX1_54 ( .A(_0__20_), .Y(_185_) );
	NOR2X1 NOR2X1_59 ( .A(_185_), .B(_182_), .Y(_186_) );
	OR2X2 OR2X2_13 ( .A(_186_), .B(_184_), .Y(_187_) );
	NOR2X1 NOR2X1_60 ( .A(b32_mode_1_bF_buf1), .B(_178_), .Y(_188_) );
	AOI22X1 AOI22X1_29 ( .A(b32_D[21]), .B(_183_), .C(_188_), .D(_187_), .Y(_189_) );
	NOR2X1 NOR2X1_61 ( .A(_184_), .B(_186_), .Y(_190_) );
	AOI21X1 AOI21X1_25 ( .A(_190_), .B(_178_), .C(_175_), .Y(_191_) );
	AOI22X1 AOI22X1_30 ( .A(_182_), .B(_175_), .C(_191_), .D(_189_), .Y(_172__1_) );
	INVX2 INVX2_5 ( .A(_0__22_), .Y(_192_) );
	NOR2X1 NOR2X1_62 ( .A(b32_mode_0_bF_buf1), .B(_179_), .Y(_193_) );
	NAND3X1 NAND3X1_9 ( .A(_0__20_), .B(_0__21_), .C(_0__22_), .Y(_194_) );
	INVX1 INVX1_55 ( .A(_194_), .Y(_195_) );
	AOI21X1 AOI21X1_26 ( .A(_0__20_), .B(_0__21_), .C(_0__22_), .Y(_196_) );
	OR2X2 OR2X2_14 ( .A(_195_), .B(_196_), .Y(_197_) );
	INVX1 INVX1_56 ( .A(b32_D[22]), .Y(_198_) );
	OAI21X1 OAI21X1_37 ( .A(_198_), .B(_177_), .C(_174_), .Y(_199_) );
	AOI21X1 AOI21X1_27 ( .A(_197_), .B(_193_), .C(_199_), .Y(_200_) );
	NOR2X1 NOR2X1_63 ( .A(b32_mode_0_bF_buf0), .B(b32_mode_1_bF_buf0), .Y(_201_) );
	NOR2X1 NOR2X1_64 ( .A(_196_), .B(_195_), .Y(_202_) );
	NAND2X1 NAND2X1_22 ( .A(_192_), .B(_184_), .Y(_203_) );
	OAI21X1 OAI21X1_38 ( .A(_0__20_), .B(_0__21_), .C(_0__22_), .Y(_204_) );
	NAND2X1 NAND2X1_23 ( .A(_204_), .B(_203_), .Y(_205_) );
	AOI22X1 AOI22X1_31 ( .A(_205_), .B(_188_), .C(_201_), .D(_202_), .Y(_206_) );
	AOI22X1 AOI22X1_32 ( .A(_192_), .B(_175_), .C(_206_), .D(_200_), .Y(_172__2_) );
	INVX4 INVX4_10 ( .A(_0__23_), .Y(_207_) );
	NOR2X1 NOR2X1_65 ( .A(_207_), .B(_194_), .Y(_208_) );
	INVX1 INVX1_57 ( .A(_208_), .Y(_209_) );
	INVX1 INVX1_58 ( .A(_201_), .Y(_210_) );
	AOI21X1 AOI21X1_28 ( .A(_207_), .B(_194_), .C(_210_), .Y(_211_) );
	INVX1 INVX1_59 ( .A(b32_D[23]), .Y(_212_) );
	OAI21X1 OAI21X1_39 ( .A(_212_), .B(_177_), .C(_174_), .Y(_213_) );
	AOI21X1 AOI21X1_29 ( .A(_209_), .B(_211_), .C(_213_), .Y(_214_) );
	NAND3X1 NAND3X1_10 ( .A(_192_), .B(_207_), .C(_184_), .Y(_215_) );
	OR2X2 OR2X2_15 ( .A(_0__20_), .B(_0__21_), .Y(_216_) );
	OAI21X1 OAI21X1_40 ( .A(_0__22_), .B(_216_), .C(_0__23_), .Y(_217_) );
	NAND2X1 NAND2X1_24 ( .A(_215_), .B(_217_), .Y(_218_) );
	XNOR2X1 XNOR2X1_5 ( .A(_196_), .B(_207_), .Y(_219_) );
	AOI22X1 AOI22X1_33 ( .A(_193_), .B(_219_), .C(_188_), .D(_218_), .Y(_220_) );
	AOI22X1 AOI22X1_34 ( .A(_207_), .B(_175_), .C(_214_), .D(_220_), .Y(_172__3_) );
	NOR2X1 NOR2X1_66 ( .A(_185_), .B(_175_), .Y(_169__0_) );
	NOR2X1 NOR2X1_67 ( .A(_182_), .B(_175_), .Y(_169__1_) );
	NOR2X1 NOR2X1_68 ( .A(_192_), .B(_175_), .Y(_169__2_) );
	NOR2X1 NOR2X1_69 ( .A(_207_), .B(_175_), .Y(_169__3_) );
	INVX1 INVX1_60 ( .A(_215_), .Y(_221_) );
	NAND2X1 NAND2X1_25 ( .A(_188_), .B(_221_), .Y(_222_) );
	AND2X2 AND2X2_5 ( .A(_196_), .B(_207_), .Y(_223_) );
	AOI22X1 AOI22X1_35 ( .A(_201_), .B(_208_), .C(_193_), .D(_223_), .Y(_224_) );
	AOI21X1 AOI21X1_30 ( .A(_222_), .B(_224_), .C(_175_), .Y(_171_) );
	NOR2X1 NOR2X1_70 ( .A(_177_), .B(_175_), .Y(_170_) );
	DFFPOSX1 DFFPOSX1_42 ( .CLK(b32_clk_bF_buf6), .D(_170_), .Q(counter_20b23_b4_load) );
	DFFPOSX1 DFFPOSX1_43 ( .CLK(b32_clk_bF_buf5), .D(_171_), .Q(counter_20b23_b4_rco) );
	DFFPOSX1 DFFPOSX1_44 ( .CLK(b32_clk_bF_buf4), .D(_169__0_), .Q(_0__20_) );
	DFFPOSX1 DFFPOSX1_45 ( .CLK(b32_clk_bF_buf3), .D(_169__1_), .Q(_0__21_) );
	DFFPOSX1 DFFPOSX1_46 ( .CLK(b32_clk_bF_buf2), .D(_169__2_), .Q(_0__22_) );
	DFFPOSX1 DFFPOSX1_47 ( .CLK(b32_clk_bF_buf1), .D(_169__3_), .Q(_0__23_) );
	DFFPOSX1 DFFPOSX1_48 ( .CLK(b32_clk_bF_buf0), .D(_172__0_), .Q(_0__20_) );
	DFFPOSX1 DFFPOSX1_49 ( .CLK(b32_clk_bF_buf7), .D(_172__1_), .Q(_0__21_) );
	DFFPOSX1 DFFPOSX1_50 ( .CLK(b32_clk_bF_buf6), .D(_172__2_), .Q(_0__22_) );
	DFFPOSX1 DFFPOSX1_51 ( .CLK(b32_clk_bF_buf5), .D(_172__3_), .Q(_0__23_) );
	INVX1 INVX1_61 ( .A(b32_enable), .Y(_229_) );
	NOR2X1 NOR2X1_71 ( .A(b32_reset), .B(_229_), .Y(_230_) );
	INVX4 INVX4_11 ( .A(_230_), .Y(_231_) );
	OAI21X1 OAI21X1_41 ( .A(b32_reset), .B(_229_), .C(_0__24_), .Y(_232_) );
	NAND2X1 NAND2X1_26 ( .A(b32_mode_0_bF_buf4), .B(b32_mode_1_bF_buf4), .Y(_233_) );
	INVX1 INVX1_62 ( .A(b32_mode_0_bF_buf3), .Y(_234_) );
	INVX1 INVX1_63 ( .A(b32_mode_1_bF_buf3), .Y(_235_) );
	OAI21X1 OAI21X1_42 ( .A(_234_), .B(_235_), .C(_0__24_), .Y(_236_) );
	OAI21X1 OAI21X1_43 ( .A(b32_D[24]), .B(_233_), .C(_236_), .Y(_237_) );
	OAI21X1 OAI21X1_44 ( .A(_231_), .B(_237_), .C(_232_), .Y(_228__0_) );
	INVX1 INVX1_64 ( .A(_0__25_), .Y(_238_) );
	INVX1 INVX1_65 ( .A(_233_), .Y(_239_) );
	NOR2X1 NOR2X1_72 ( .A(_0__24_), .B(_0__25_), .Y(_240_) );
	INVX1 INVX1_66 ( .A(_0__24_), .Y(_241_) );
	NOR2X1 NOR2X1_73 ( .A(_241_), .B(_238_), .Y(_242_) );
	OR2X2 OR2X2_16 ( .A(_242_), .B(_240_), .Y(_243_) );
	NOR2X1 NOR2X1_74 ( .A(b32_mode_1_bF_buf2), .B(_234_), .Y(_244_) );
	AOI22X1 AOI22X1_36 ( .A(b32_D[25]), .B(_239_), .C(_244_), .D(_243_), .Y(_245_) );
	NOR2X1 NOR2X1_75 ( .A(_240_), .B(_242_), .Y(_246_) );
	AOI21X1 AOI21X1_31 ( .A(_246_), .B(_234_), .C(_231_), .Y(_247_) );
	AOI22X1 AOI22X1_37 ( .A(_238_), .B(_231_), .C(_247_), .D(_245_), .Y(_228__1_) );
	INVX2 INVX2_6 ( .A(_0__26_), .Y(_248_) );
	NOR2X1 NOR2X1_76 ( .A(b32_mode_0_bF_buf2), .B(_235_), .Y(_249_) );
	NAND3X1 NAND3X1_11 ( .A(_0__24_), .B(_0__25_), .C(_0__26_), .Y(_250_) );
	INVX1 INVX1_67 ( .A(_250_), .Y(_251_) );
	AOI21X1 AOI21X1_32 ( .A(_0__24_), .B(_0__25_), .C(_0__26_), .Y(_252_) );
	OR2X2 OR2X2_17 ( .A(_251_), .B(_252_), .Y(_253_) );
	INVX1 INVX1_68 ( .A(b32_D[26]), .Y(_254_) );
	OAI21X1 OAI21X1_45 ( .A(_254_), .B(_233_), .C(_230_), .Y(_255_) );
	AOI21X1 AOI21X1_33 ( .A(_253_), .B(_249_), .C(_255_), .Y(_256_) );
	NOR2X1 NOR2X1_77 ( .A(b32_mode_0_bF_buf1), .B(b32_mode_1_bF_buf1), .Y(_257_) );
	NOR2X1 NOR2X1_78 ( .A(_252_), .B(_251_), .Y(_258_) );
	NAND2X1 NAND2X1_27 ( .A(_248_), .B(_240_), .Y(_259_) );
	OAI21X1 OAI21X1_46 ( .A(_0__24_), .B(_0__25_), .C(_0__26_), .Y(_260_) );
	NAND2X1 NAND2X1_28 ( .A(_260_), .B(_259_), .Y(_261_) );
	AOI22X1 AOI22X1_38 ( .A(_261_), .B(_244_), .C(_257_), .D(_258_), .Y(_262_) );
	AOI22X1 AOI22X1_39 ( .A(_248_), .B(_231_), .C(_262_), .D(_256_), .Y(_228__2_) );
	INVX4 INVX4_12 ( .A(_0__27_), .Y(_263_) );
	NOR2X1 NOR2X1_79 ( .A(_263_), .B(_250_), .Y(_264_) );
	INVX1 INVX1_69 ( .A(_264_), .Y(_265_) );
	INVX1 INVX1_70 ( .A(_257_), .Y(_266_) );
	AOI21X1 AOI21X1_34 ( .A(_263_), .B(_250_), .C(_266_), .Y(_267_) );
	INVX1 INVX1_71 ( .A(b32_D[27]), .Y(_268_) );
	OAI21X1 OAI21X1_47 ( .A(_268_), .B(_233_), .C(_230_), .Y(_269_) );
	AOI21X1 AOI21X1_35 ( .A(_265_), .B(_267_), .C(_269_), .Y(_270_) );
	NAND3X1 NAND3X1_12 ( .A(_248_), .B(_263_), .C(_240_), .Y(_271_) );
	OR2X2 OR2X2_18 ( .A(_0__24_), .B(_0__25_), .Y(_272_) );
	OAI21X1 OAI21X1_48 ( .A(_0__26_), .B(_272_), .C(_0__27_), .Y(_273_) );
	NAND2X1 NAND2X1_29 ( .A(_271_), .B(_273_), .Y(_274_) );
	XNOR2X1 XNOR2X1_6 ( .A(_252_), .B(_263_), .Y(_275_) );
	AOI22X1 AOI22X1_40 ( .A(_249_), .B(_275_), .C(_244_), .D(_274_), .Y(_276_) );
	AOI22X1 AOI22X1_41 ( .A(_263_), .B(_231_), .C(_270_), .D(_276_), .Y(_228__3_) );
	NOR2X1 NOR2X1_80 ( .A(_241_), .B(_231_), .Y(_225__0_) );
	NOR2X1 NOR2X1_81 ( .A(_238_), .B(_231_), .Y(_225__1_) );
	NOR2X1 NOR2X1_82 ( .A(_248_), .B(_231_), .Y(_225__2_) );
	NOR2X1 NOR2X1_83 ( .A(_263_), .B(_231_), .Y(_225__3_) );
	INVX1 INVX1_72 ( .A(_271_), .Y(_277_) );
	NAND2X1 NAND2X1_30 ( .A(_244_), .B(_277_), .Y(_278_) );
	AND2X2 AND2X2_6 ( .A(_252_), .B(_263_), .Y(_279_) );
	AOI22X1 AOI22X1_42 ( .A(_257_), .B(_264_), .C(_249_), .D(_279_), .Y(_280_) );
	AOI21X1 AOI21X1_36 ( .A(_278_), .B(_280_), .C(_231_), .Y(_227_) );
	NOR2X1 NOR2X1_84 ( .A(_233_), .B(_231_), .Y(_226_) );
	DFFPOSX1 DFFPOSX1_52 ( .CLK(b32_clk_bF_buf4), .D(_226_), .Q(counter_24b27_b4_load) );
	DFFPOSX1 DFFPOSX1_53 ( .CLK(b32_clk_bF_buf3), .D(_227_), .Q(counter_24b27_b4_rco) );
	DFFPOSX1 DFFPOSX1_54 ( .CLK(b32_clk_bF_buf2), .D(_225__0_), .Q(_0__24_) );
	DFFPOSX1 DFFPOSX1_55 ( .CLK(b32_clk_bF_buf1), .D(_225__1_), .Q(_0__25_) );
	DFFPOSX1 DFFPOSX1_56 ( .CLK(b32_clk_bF_buf0), .D(_225__2_), .Q(_0__26_) );
	DFFPOSX1 DFFPOSX1_57 ( .CLK(b32_clk_bF_buf7), .D(_225__3_), .Q(_0__27_) );
	DFFPOSX1 DFFPOSX1_58 ( .CLK(b32_clk_bF_buf6), .D(_228__0_), .Q(_0__24_) );
	DFFPOSX1 DFFPOSX1_59 ( .CLK(b32_clk_bF_buf5), .D(_228__1_), .Q(_0__25_) );
	DFFPOSX1 DFFPOSX1_60 ( .CLK(b32_clk_bF_buf4), .D(_228__2_), .Q(_0__26_) );
	DFFPOSX1 DFFPOSX1_61 ( .CLK(b32_clk_bF_buf3), .D(_228__3_), .Q(_0__27_) );
	INVX1 INVX1_73 ( .A(b32_enable), .Y(_285_) );
	NOR2X1 NOR2X1_85 ( .A(b32_reset), .B(_285_), .Y(_286_) );
	INVX4 INVX4_13 ( .A(_286_), .Y(_287_) );
	OAI21X1 OAI21X1_49 ( .A(b32_reset), .B(_285_), .C(_0__28_), .Y(_288_) );
	NAND2X1 NAND2X1_31 ( .A(b32_mode_0_bF_buf0), .B(b32_mode_1_bF_buf0), .Y(_289_) );
	INVX1 INVX1_74 ( .A(b32_mode_0_bF_buf4), .Y(_290_) );
	INVX1 INVX1_75 ( .A(b32_mode_1_bF_buf4), .Y(_291_) );
	OAI21X1 OAI21X1_50 ( .A(_290_), .B(_291_), .C(_0__28_), .Y(_292_) );
	OAI21X1 OAI21X1_51 ( .A(b32_D[28]), .B(_289_), .C(_292_), .Y(_293_) );
	OAI21X1 OAI21X1_52 ( .A(_287_), .B(_293_), .C(_288_), .Y(_284__0_) );
	INVX1 INVX1_76 ( .A(_0__29_), .Y(_294_) );
	INVX1 INVX1_77 ( .A(_289_), .Y(_295_) );
	NOR2X1 NOR2X1_86 ( .A(_0__28_), .B(_0__29_), .Y(_296_) );
	INVX1 INVX1_78 ( .A(_0__28_), .Y(_297_) );
	NOR2X1 NOR2X1_87 ( .A(_297_), .B(_294_), .Y(_298_) );
	OR2X2 OR2X2_19 ( .A(_298_), .B(_296_), .Y(_299_) );
	NOR2X1 NOR2X1_88 ( .A(b32_mode_1_bF_buf3), .B(_290_), .Y(_300_) );
	AOI22X1 AOI22X1_43 ( .A(b32_D[29]), .B(_295_), .C(_300_), .D(_299_), .Y(_301_) );
	NOR2X1 NOR2X1_89 ( .A(_296_), .B(_298_), .Y(_302_) );
	AOI21X1 AOI21X1_37 ( .A(_302_), .B(_290_), .C(_287_), .Y(_303_) );
	AOI22X1 AOI22X1_44 ( .A(_294_), .B(_287_), .C(_303_), .D(_301_), .Y(_284__1_) );
	INVX2 INVX2_7 ( .A(_0__30_), .Y(_304_) );
	NOR2X1 NOR2X1_90 ( .A(b32_mode_0_bF_buf3), .B(_291_), .Y(_305_) );
	NAND3X1 NAND3X1_13 ( .A(_0__28_), .B(_0__29_), .C(_0__30_), .Y(_306_) );
	INVX1 INVX1_79 ( .A(_306_), .Y(_307_) );
	AOI21X1 AOI21X1_38 ( .A(_0__28_), .B(_0__29_), .C(_0__30_), .Y(_308_) );
	OR2X2 OR2X2_20 ( .A(_307_), .B(_308_), .Y(_309_) );
	INVX1 INVX1_80 ( .A(b32_D[30]), .Y(_310_) );
	OAI21X1 OAI21X1_53 ( .A(_310_), .B(_289_), .C(_286_), .Y(_311_) );
	AOI21X1 AOI21X1_39 ( .A(_309_), .B(_305_), .C(_311_), .Y(_312_) );
	NOR2X1 NOR2X1_91 ( .A(b32_mode_0_bF_buf2), .B(b32_mode_1_bF_buf2), .Y(_313_) );
	NOR2X1 NOR2X1_92 ( .A(_308_), .B(_307_), .Y(_314_) );
	NAND2X1 NAND2X1_32 ( .A(_304_), .B(_296_), .Y(_315_) );
	OAI21X1 OAI21X1_54 ( .A(_0__28_), .B(_0__29_), .C(_0__30_), .Y(_316_) );
	NAND2X1 NAND2X1_33 ( .A(_316_), .B(_315_), .Y(_317_) );
	AOI22X1 AOI22X1_45 ( .A(_317_), .B(_300_), .C(_313_), .D(_314_), .Y(_318_) );
	AOI22X1 AOI22X1_46 ( .A(_304_), .B(_287_), .C(_318_), .D(_312_), .Y(_284__2_) );
	INVX4 INVX4_14 ( .A(_0__31_), .Y(_319_) );
	NOR2X1 NOR2X1_93 ( .A(_319_), .B(_306_), .Y(_320_) );
	INVX1 INVX1_81 ( .A(_320_), .Y(_321_) );
	INVX1 INVX1_82 ( .A(_313_), .Y(_322_) );
	AOI21X1 AOI21X1_40 ( .A(_319_), .B(_306_), .C(_322_), .Y(_323_) );
	INVX1 INVX1_83 ( .A(b32_D[31]), .Y(_324_) );
	OAI21X1 OAI21X1_55 ( .A(_324_), .B(_289_), .C(_286_), .Y(_325_) );
	AOI21X1 AOI21X1_41 ( .A(_321_), .B(_323_), .C(_325_), .Y(_326_) );
	NAND3X1 NAND3X1_14 ( .A(_304_), .B(_319_), .C(_296_), .Y(_327_) );
	OR2X2 OR2X2_21 ( .A(_0__28_), .B(_0__29_), .Y(_328_) );
	OAI21X1 OAI21X1_56 ( .A(_0__30_), .B(_328_), .C(_0__31_), .Y(_329_) );
	NAND2X1 NAND2X1_34 ( .A(_327_), .B(_329_), .Y(_330_) );
	XNOR2X1 XNOR2X1_7 ( .A(_308_), .B(_319_), .Y(_331_) );
	AOI22X1 AOI22X1_47 ( .A(_305_), .B(_331_), .C(_300_), .D(_330_), .Y(_332_) );
	AOI22X1 AOI22X1_48 ( .A(_319_), .B(_287_), .C(_326_), .D(_332_), .Y(_284__3_) );
	NOR2X1 NOR2X1_94 ( .A(_297_), .B(_287_), .Y(_281__0_) );
	NOR2X1 NOR2X1_95 ( .A(_294_), .B(_287_), .Y(_281__1_) );
	NOR2X1 NOR2X1_96 ( .A(_304_), .B(_287_), .Y(_281__2_) );
	NOR2X1 NOR2X1_97 ( .A(_319_), .B(_287_), .Y(_281__3_) );
	INVX1 INVX1_84 ( .A(_327_), .Y(_333_) );
	NAND2X1 NAND2X1_35 ( .A(_300_), .B(_333_), .Y(_334_) );
	AND2X2 AND2X2_7 ( .A(_308_), .B(_319_), .Y(_335_) );
	AOI22X1 AOI22X1_49 ( .A(_313_), .B(_320_), .C(_305_), .D(_335_), .Y(_336_) );
	AOI21X1 AOI21X1_42 ( .A(_334_), .B(_336_), .C(_287_), .Y(_283_) );
	NOR2X1 NOR2X1_98 ( .A(_289_), .B(_287_), .Y(_282_) );
	DFFPOSX1 DFFPOSX1_62 ( .CLK(b32_clk_bF_buf2), .D(_282_), .Q(counter_28b31_b4_load) );
	DFFPOSX1 DFFPOSX1_63 ( .CLK(b32_clk_bF_buf1), .D(_283_), .Q(counter_28b31_b4_rco) );
	DFFPOSX1 DFFPOSX1_64 ( .CLK(b32_clk_bF_buf0), .D(_281__0_), .Q(_0__28_) );
	DFFPOSX1 DFFPOSX1_65 ( .CLK(b32_clk_bF_buf7), .D(_281__1_), .Q(_0__29_) );
	DFFPOSX1 DFFPOSX1_66 ( .CLK(b32_clk_bF_buf6), .D(_281__2_), .Q(_0__30_) );
	DFFPOSX1 DFFPOSX1_67 ( .CLK(b32_clk_bF_buf5), .D(_281__3_), .Q(_0__31_) );
	DFFPOSX1 DFFPOSX1_68 ( .CLK(b32_clk_bF_buf4), .D(_284__0_), .Q(_0__28_) );
	DFFPOSX1 DFFPOSX1_69 ( .CLK(b32_clk_bF_buf3), .D(_284__1_), .Q(_0__29_) );
	DFFPOSX1 DFFPOSX1_70 ( .CLK(b32_clk_bF_buf2), .D(_284__2_), .Q(_0__30_) );
	DFFPOSX1 DFFPOSX1_71 ( .CLK(b32_clk_bF_buf1), .D(_284__3_), .Q(_0__31_) );
	INVX1 INVX1_85 ( .A(b32_enable), .Y(_341_) );
	NOR2X1 NOR2X1_99 ( .A(b32_reset), .B(_341_), .Y(_342_) );
	INVX4 INVX4_15 ( .A(_342_), .Y(_343_) );
	OAI21X1 OAI21X1_57 ( .A(b32_reset), .B(_341_), .C(_0__4_), .Y(_344_) );
	NAND2X1 NAND2X1_36 ( .A(b32_mode_0_bF_buf1), .B(b32_mode_1_bF_buf1), .Y(_345_) );
	INVX1 INVX1_86 ( .A(b32_mode_0_bF_buf0), .Y(_346_) );
	INVX1 INVX1_87 ( .A(b32_mode_1_bF_buf0), .Y(_347_) );
	OAI21X1 OAI21X1_58 ( .A(_346_), .B(_347_), .C(_0__4_), .Y(_348_) );
	OAI21X1 OAI21X1_59 ( .A(b32_D[4]), .B(_345_), .C(_348_), .Y(_349_) );
	OAI21X1 OAI21X1_60 ( .A(_343_), .B(_349_), .C(_344_), .Y(_340__0_) );
	INVX1 INVX1_88 ( .A(_0__5_), .Y(_350_) );
	INVX1 INVX1_89 ( .A(_345_), .Y(_351_) );
	NOR2X1 NOR2X1_100 ( .A(_0__4_), .B(_0__5_), .Y(_352_) );
	INVX1 INVX1_90 ( .A(_0__4_), .Y(_353_) );
	NOR2X1 NOR2X1_101 ( .A(_353_), .B(_350_), .Y(_354_) );
	OR2X2 OR2X2_22 ( .A(_354_), .B(_352_), .Y(_355_) );
	NOR2X1 NOR2X1_102 ( .A(b32_mode_1_bF_buf4), .B(_346_), .Y(_356_) );
	AOI22X1 AOI22X1_50 ( .A(b32_D[5]), .B(_351_), .C(_356_), .D(_355_), .Y(_357_) );
	NOR2X1 NOR2X1_103 ( .A(_352_), .B(_354_), .Y(_358_) );
	AOI21X1 AOI21X1_43 ( .A(_358_), .B(_346_), .C(_343_), .Y(_359_) );
	AOI22X1 AOI22X1_51 ( .A(_350_), .B(_343_), .C(_359_), .D(_357_), .Y(_340__1_) );
	INVX2 INVX2_8 ( .A(_0__6_), .Y(_360_) );
	NOR2X1 NOR2X1_104 ( .A(b32_mode_0_bF_buf4), .B(_347_), .Y(_361_) );
	NAND3X1 NAND3X1_15 ( .A(_0__4_), .B(_0__5_), .C(_0__6_), .Y(_362_) );
	INVX1 INVX1_91 ( .A(_362_), .Y(_363_) );
	AOI21X1 AOI21X1_44 ( .A(_0__4_), .B(_0__5_), .C(_0__6_), .Y(_364_) );
	OR2X2 OR2X2_23 ( .A(_363_), .B(_364_), .Y(_365_) );
	INVX1 INVX1_92 ( .A(b32_D[6]), .Y(_366_) );
	OAI21X1 OAI21X1_61 ( .A(_366_), .B(_345_), .C(_342_), .Y(_367_) );
	AOI21X1 AOI21X1_45 ( .A(_365_), .B(_361_), .C(_367_), .Y(_368_) );
	NOR2X1 NOR2X1_105 ( .A(b32_mode_0_bF_buf3), .B(b32_mode_1_bF_buf3), .Y(_369_) );
	NOR2X1 NOR2X1_106 ( .A(_364_), .B(_363_), .Y(_370_) );
	NAND2X1 NAND2X1_37 ( .A(_360_), .B(_352_), .Y(_371_) );
	OAI21X1 OAI21X1_62 ( .A(_0__4_), .B(_0__5_), .C(_0__6_), .Y(_372_) );
	NAND2X1 NAND2X1_38 ( .A(_372_), .B(_371_), .Y(_373_) );
	AOI22X1 AOI22X1_52 ( .A(_373_), .B(_356_), .C(_369_), .D(_370_), .Y(_374_) );
	AOI22X1 AOI22X1_53 ( .A(_360_), .B(_343_), .C(_374_), .D(_368_), .Y(_340__2_) );
	INVX4 INVX4_16 ( .A(_0__7_), .Y(_375_) );
	NOR2X1 NOR2X1_107 ( .A(_375_), .B(_362_), .Y(_376_) );
	INVX1 INVX1_93 ( .A(_376_), .Y(_377_) );
	INVX1 INVX1_94 ( .A(_369_), .Y(_378_) );
	AOI21X1 AOI21X1_46 ( .A(_375_), .B(_362_), .C(_378_), .Y(_379_) );
	INVX1 INVX1_95 ( .A(b32_D[7]), .Y(_380_) );
	OAI21X1 OAI21X1_63 ( .A(_380_), .B(_345_), .C(_342_), .Y(_381_) );
	AOI21X1 AOI21X1_47 ( .A(_377_), .B(_379_), .C(_381_), .Y(_382_) );
	NAND3X1 NAND3X1_16 ( .A(_360_), .B(_375_), .C(_352_), .Y(_383_) );
	OR2X2 OR2X2_24 ( .A(_0__4_), .B(_0__5_), .Y(_384_) );
	OAI21X1 OAI21X1_64 ( .A(_0__6_), .B(_384_), .C(_0__7_), .Y(_385_) );
	NAND2X1 NAND2X1_39 ( .A(_383_), .B(_385_), .Y(_386_) );
	XNOR2X1 XNOR2X1_8 ( .A(_364_), .B(_375_), .Y(_387_) );
	AOI22X1 AOI22X1_54 ( .A(_361_), .B(_387_), .C(_356_), .D(_386_), .Y(_388_) );
	AOI22X1 AOI22X1_55 ( .A(_375_), .B(_343_), .C(_382_), .D(_388_), .Y(_340__3_) );
	NOR2X1 NOR2X1_108 ( .A(_353_), .B(_343_), .Y(_337__0_) );
	NOR2X1 NOR2X1_109 ( .A(_350_), .B(_343_), .Y(_337__1_) );
	NOR2X1 NOR2X1_110 ( .A(_360_), .B(_343_), .Y(_337__2_) );
	NOR2X1 NOR2X1_111 ( .A(_375_), .B(_343_), .Y(_337__3_) );
	INVX1 INVX1_96 ( .A(_383_), .Y(_389_) );
	NAND2X1 NAND2X1_40 ( .A(_356_), .B(_389_), .Y(_390_) );
	AND2X2 AND2X2_8 ( .A(_364_), .B(_375_), .Y(_391_) );
	AOI22X1 AOI22X1_56 ( .A(_369_), .B(_376_), .C(_361_), .D(_391_), .Y(_392_) );
	AOI21X1 AOI21X1_48 ( .A(_390_), .B(_392_), .C(_343_), .Y(_339_) );
	NOR2X1 NOR2X1_112 ( .A(_345_), .B(_343_), .Y(_338_) );
	DFFPOSX1 DFFPOSX1_72 ( .CLK(b32_clk_bF_buf0), .D(_338_), .Q(counter_4b7_b4_load) );
	DFFPOSX1 DFFPOSX1_73 ( .CLK(b32_clk_bF_buf7), .D(_339_), .Q(counter_4b7_b4_rco) );
	DFFPOSX1 DFFPOSX1_74 ( .CLK(b32_clk_bF_buf6), .D(_337__0_), .Q(_0__4_) );
	DFFPOSX1 DFFPOSX1_75 ( .CLK(b32_clk_bF_buf5), .D(_337__1_), .Q(_0__5_) );
	DFFPOSX1 DFFPOSX1_76 ( .CLK(b32_clk_bF_buf4), .D(_337__2_), .Q(_0__6_) );
	DFFPOSX1 DFFPOSX1_77 ( .CLK(b32_clk_bF_buf3), .D(_337__3_), .Q(_0__7_) );
	DFFPOSX1 DFFPOSX1_78 ( .CLK(b32_clk_bF_buf2), .D(_340__0_), .Q(_0__4_) );
	DFFPOSX1 DFFPOSX1_79 ( .CLK(b32_clk_bF_buf1), .D(_340__1_), .Q(_0__5_) );
	DFFPOSX1 DFFPOSX1_80 ( .CLK(b32_clk_bF_buf0), .D(_340__2_), .Q(_0__6_) );
endmodule
