*** SPICE deck for cell AOI22{lay} from library Design_NOR3_NAND3_AOI22
*** Created on Sun Dec 06, 2020 17:40:10
*** Last revised on Sun Dec 06, 2020 18:08:08
*** Written on Sun Dec 06, 2020 18:45:20 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

*** TOP LEVEL CELL: AOI22{lay}
Mnmos@0 OUT A_or_B GND GND_or NMOS L=0.2U W=0.3U AS=1.28P AD=0.353P PS=7.2U PD=2.4U
Mnmos@1 GND_or A_and_B_0 A_or_B GND_or NMOS L=0.2U W=0.3U AS=0.487P AD=0.405P PS=2.867U PD=2.7U
Mnmos@2 A_or_B A GND_or GND_or NMOS L=0.2U W=0.3U AS=0.405P AD=0.487P PS=2.7U PD=2.867U
Mnmos@3 A B_1 net@52 GND_or NMOS L=0.2U W=0.6U AS=0.128P AD=0.307P PS=1.05U PD=1.8U
Mnmos@4 net@52 A_1 GND_AND1 GND_or NMOS L=0.2U W=0.6U AS=1.36P AD=0.128P PS=7.4U PD=1.05U
Mnmos@5 A_and_B_0 B_0 net@75 GND_or NMOS L=0.2U W=0.6U AS=0.128P AD=0.307P PS=1.05U PD=1.8U
Mnmos@6 net@75 A_0 GND_AND0 GND_or NMOS L=0.2U W=0.6U AS=1.36P AD=0.128P PS=7.4U PD=1.05U
Mpmos@0 VDD A_or_B OUT VDD_or PMOS L=0.2U W=0.7U AS=0.353P AD=1.42P PS=2.4U PD=7.6U
Mpmos@1 A_or_B A_and_B_0 net@36 VDD_or PMOS L=0.2U W=1.5U AS=0.375P AD=0.487P PS=2U PD=2.867U
Mpmos@2 net@36 A VDD_or VDD_or PMOS L=0.2U W=1.5U AS=1.4P AD=0.375P PS=7.2U PD=2U
Mpmos@3 VDD_AND1 A_1 A VDD_or PMOS L=0.2U W=0.8U AS=0.307P AD=1.105P PS=1.8U PD=5.8U
Mpmos@4 A B_1 VDD_AND1 VDD_or PMOS L=0.2U W=0.8U AS=1.105P AD=0.307P PS=5.8U PD=1.8U
Mpmos@5 VDD_AND0 A_0 A_and_B_0 VDD_or PMOS L=0.2U W=0.8U AS=0.307P AD=1.105P PS=1.8U PD=5.8U
Mpmos@6 A_and_B_0 B_0 VDD_AND0 VDD_or PMOS L=0.2U W=0.8U AS=1.105P AD=0.307P PS=5.8U PD=1.8U
.END
