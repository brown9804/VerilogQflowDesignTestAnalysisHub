*** SPICE deck for cell NOR3{lay} from library Design_NOR3_NAND3_AOI22
*** Created on Sun Dec 06, 2020 18:26:05
*** Last revised on Sun Dec 06, 2020 18:43:16
*** Written on Sun Dec 06, 2020 18:44:54 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

*** TOP LEVEL CELL: NOR3{lay}
Mnmos@3 X_or_W_or_Z X gnd gnd NMOS L=0.2U W=0.3U AS=0.973P AD=0.459P PS=5.017U PD=2.575U
Mnmos@4 gnd W X_or_W_or_Z gnd NMOS L=0.2U W=0.3U AS=0.459P AD=0.973P PS=2.575U PD=5.017U
Mnmos@5 X_or_W_or_Z Z gnd gnd NMOS L=0.2U W=0.3U AS=0.973P AD=0.459P PS=5.017U PD=2.575U
Mpmos@3 vdd X net@60 vdd PMOS L=0.2U W=1.9U AS=0.57P AD=2.94P PS=2.5U PD=13.2U
Mpmos@4 net@60 W net@61 vdd PMOS L=0.2U W=1.9U AS=0.57P AD=0.57P PS=2.5U PD=2.5U
Mpmos@5 net@61 Z X_or_W_or_Z vdd PMOS L=0.2U W=1.9U AS=0.459P AD=0.57P PS=2.575U PD=2.5U
.END
