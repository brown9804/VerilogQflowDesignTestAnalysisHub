module uart ( gnd, vdd, reset, txclk, ld_tx_data, tx_data, tx_enable, rxclk, uld_rx_data, rx_enable, rx_in, tx_out, tx_empty, rx_data, rx_empty);

input gnd, vdd;
input reset;
input txclk;
input ld_tx_data;
input tx_enable;
input rxclk;
input uld_rx_data;
input rx_enable;
input rx_in;
output tx_out;
output tx_empty;
output rx_empty;
input [7:0] tx_data;
output [7:0] rx_data;

	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(rxclk), .Y(rxclk_bF_buf4) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(rxclk), .Y(rxclk_bF_buf3) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(rxclk), .Y(rxclk_bF_buf2) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(rxclk), .Y(rxclk_bF_buf1) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(rxclk), .Y(rxclk_bF_buf0) );
	BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_162_), .Y(_162__bF_buf5) );
	BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_162_), .Y(_162__bF_buf4) );
	BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_162_), .Y(_162__bF_buf3) );
	BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_162_), .Y(_162__bF_buf2) );
	BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_162_), .Y(_162__bF_buf1) );
	BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(_162_), .Y(_162__bF_buf0) );
	BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data), .Y(uld_rx_data_bF_buf3) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data), .Y(uld_rx_data_bF_buf2) );
	BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data), .Y(uld_rx_data_bF_buf1) );
	BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data), .Y(uld_rx_data_bF_buf0) );
	INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(rx_d2), .Y(_163_) );
	INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_0_), .Y(_164_) );
	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_1_), .B(_164_), .Y(_165_) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_3_), .Y(_166_) );
	INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_2_), .Y(_10_) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_1_), .B(rx_cnt_0_), .Y(_11_) );
	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_11_), .Y(_12_) );
	XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_166_), .Y(_13_) );
	OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_1_), .B(rx_cnt_0_), .C(rx_cnt_2_), .Y(_14_) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_12_), .Y(_15_) );
	INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(rx_enable), .Y(_16_) );
	NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(rx_sample_cnt_1_), .B(rx_sample_cnt_0_), .C(rx_sample_cnt_2_), .Y(_17_) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(rx_sample_cnt_3_), .Y(_18_) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(rx_busy), .B(_18_), .Y(_19_) );
	NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_17_), .C(_19_), .Y(_20_) );
	AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_15_), .Y(_21_) );
	NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_13_), .C(_21_), .Y(_22_) );
	NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_4_), .B(_22_), .Y(_23_) );
	OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_22_), .C(_23_), .Y(_4__4_) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_20_), .Y(_24_) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_3_), .B(_10_), .Y(_25_) );
	NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_25_), .Y(_26_) );
	OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_26_), .Y(_27_) );
	OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_24_), .C(rx_reg_3_), .Y(_28_) );
	OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_27_), .C(_28_), .Y(_4__3_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_3_), .B(_15_), .Y(_29_) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_1_), .Y(_30_) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_164_), .Y(_31_) );
	NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_31_), .C(_29_), .Y(_32_) );
	NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_2_), .B(_32_), .Y(_33_) );
	OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_32_), .C(_33_), .Y(_4__2_) );
	NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_0_), .B(_30_), .Y(_34_) );
	NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_34_), .C(_29_), .Y(_35_) );
	NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_1_), .B(_35_), .Y(_36_) );
	OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_35_), .C(_36_), .Y(_4__1_) );
	NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_20_), .C(_29_), .Y(_37_) );
	NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_0_), .B(_37_), .Y(_38_) );
	OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_37_), .C(_38_), .Y(_4__0_) );
	OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(rx_busy), .B(_163_), .C(rx_enable), .Y(_39_) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_39_), .Y(_40_) );
	OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(rx_sample_cnt_3_), .B(_17_), .C(rx_busy), .Y(_41_) );
	AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_41_), .Y(_42_) );
	NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_3_), .B(rx_cnt_2_), .Y(_43_) );
	NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_43_), .Y(_44_) );
	OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_44_), .C(_164_), .Y(_45_) );
	OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_45_), .C(_164_), .D(_42_), .Y(_1__0_) );
	OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_34_), .C(_20_), .Y(_46_) );
	OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_42_), .C(_46_), .Y(_1__1_) );
	NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(rx_enable), .B(_31_), .Y(_47_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_47_), .Y(_48_) );
	NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_19_), .Y(_49_) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_50_) );
	AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_2_), .B(_31_), .C(_50_), .Y(_51_) );
	OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_2_), .B(_48_), .C(_51_), .Y(_52_) );
	OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_42_), .C(_52_), .Y(_1__2_) );
	NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_25_), .C(_48_), .Y(_53_) );
	INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_42_), .Y(_54_) );
	OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_54_), .C(rx_cnt_3_), .Y(_55_) );
	NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_55_), .Y(_1__3_) );
	INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(rx_sample_cnt_0_), .Y(_56_) );
	NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_16_), .Y(_57_) );
	AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(rx_busy), .C(_56_), .D(_39_), .Y(_5__0_) );
	INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(rx_sample_cnt_1_), .Y(_58_) );
	NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(rx_sample_cnt_1_), .B(rx_sample_cnt_0_), .Y(_59_) );
	AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(rx_busy), .Y(_60_) );
	OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(rx_sample_cnt_1_), .B(_57_), .C(_60_), .Y(_61_) );
	OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_40_), .C(_61_), .Y(_5__1_) );
	INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(rx_sample_cnt_2_), .Y(_62_) );
	AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(rx_busy), .Y(_63_) );
	OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_59_), .C(_62_), .Y(_64_) );
	NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_63_), .Y(_65_) );
	OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_40_), .C(_65_), .Y(_5__2_) );
	OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_63_), .C(rx_sample_cnt_3_), .Y(_66_) );
	OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_50_), .C(_66_), .Y(_5__3_) );
	NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(uld_rx_data_bF_buf3), .Y(_67_) );
	NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(rx_cnt_3_), .B(_10_), .C(_165_), .Y(_68_) );
	NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_68_), .Y(_69_) );
	AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_20_), .C(_67_), .Y(_3_) );
	INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_167__0_), .Y(_70_) );
	NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_0_), .B(uld_rx_data_bF_buf2), .Y(_71_) );
	OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf1), .B(_70_), .C(_71_), .Y(_2__0_) );
	INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_167__1_), .Y(_72_) );
	NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_1_), .B(uld_rx_data_bF_buf0), .Y(_73_) );
	OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf3), .B(_72_), .C(_73_), .Y(_2__1_) );
	INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_167__2_), .Y(_74_) );
	NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_2_), .B(uld_rx_data_bF_buf2), .Y(_75_) );
	OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf1), .B(_74_), .C(_75_), .Y(_2__2_) );
	INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_167__3_), .Y(_76_) );
	NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_3_), .B(uld_rx_data_bF_buf0), .Y(_77_) );
	OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf3), .B(_76_), .C(_77_), .Y(_2__3_) );
	INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_167__4_), .Y(_78_) );
	NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_4_), .B(uld_rx_data_bF_buf2), .Y(_79_) );
	OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf1), .B(_78_), .C(_79_), .Y(_2__4_) );
	INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_167__5_), .Y(_80_) );
	NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf0), .B(rx_reg_5_), .Y(_81_) );
	OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf3), .B(_80_), .C(_81_), .Y(_2__5_) );
	INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_6_), .Y(_82_) );
	NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf2), .B(_167__6_), .Y(_83_) );
	AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf1), .B(_82_), .C(_83_), .Y(_2__6_) );
	INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_7_), .Y(_84_) );
	NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf0), .B(_167__7_), .Y(_85_) );
	AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(uld_rx_data_bF_buf3), .B(_84_), .C(_85_), .Y(_2__7_) );
	INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_0_), .Y(_86_) );
	OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_86_), .C(tx_enable), .Y(_87_) );
	AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_169_), .C(_87_), .Y(_6__0_) );
	INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(tx_enable), .Y(_88_) );
	NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_88_), .Y(_89_) );
	NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_2_), .B(tx_cnt_1_), .Y(_90_) );
	NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_0_), .B(tx_cnt_3_), .C(_90_), .Y(_91_) );
	NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_0_), .B(tx_cnt_1_), .Y(_92_) );
	NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_0_), .B(tx_cnt_1_), .Y(_93_) );
	INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_94_) );
	NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_94_), .Y(_95_) );
	NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_91_), .C(_95_), .Y(_96_) );
	OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_88_), .C(tx_cnt_1_), .Y(_97_) );
	AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_97_), .C(_88_), .Y(_6__1_) );
	INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_2_), .Y(_98_) );
	INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_89_), .Y(_99_) );
	OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_99_), .C(_98_), .Y(_100_) );
	NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_89_), .Y(_101_) );
	OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_98_), .Y(_102_) );
	NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_102_), .Y(_103_) );
	NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_103_), .Y(_6__2_) );
	OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_91_), .C(tx_enable), .Y(_104_) );
	OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_101_), .C(tx_cnt_3_), .Y(_105_) );
	OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(tx_cnt_3_), .Y(_106_) );
	AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_105_), .C(_104_), .Y(_6__3_) );
	INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(tx_reg_0_), .Y(_107_) );
	INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(tx_data[0]), .Y(_108_) );
	AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(ld_tx_data), .Y(_109_) );
	MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_107_), .S(_109_), .Y(_9__0_) );
	INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(tx_reg_1_), .Y(_110_) );
	INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(tx_data[1]), .Y(_111_) );
	MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_110_), .S(_109_), .Y(_9__1_) );
	INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(tx_reg_2_), .Y(_112_) );
	INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(tx_data[2]), .Y(_113_) );
	MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_112_), .S(_109_), .Y(_9__2_) );
	INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(tx_reg_3_), .Y(_114_) );
	INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(tx_data[3]), .Y(_115_) );
	MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_114_), .S(_109_), .Y(_9__3_) );
	INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(tx_reg_4_), .Y(_116_) );
	INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(tx_data[4]), .Y(_117_) );
	MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_116_), .S(_109_), .Y(_9__4_) );
	INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(tx_reg_5_), .Y(_118_) );
	INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(tx_data[5]), .Y(_119_) );
	MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_118_), .S(_109_), .Y(_9__5_) );
	INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(tx_data[6]), .Y(_120_) );
	NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(tx_reg_6_), .B(_109_), .Y(_121_) );
	AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_109_), .C(_121_), .Y(_9__6_) );
	INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(tx_data[7]), .Y(_122_) );
	NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(tx_reg_7_), .B(_109_), .Y(_123_) );
	AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_109_), .C(_123_), .Y(_9__7_) );
	INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_169_), .Y(_124_) );
	OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(ld_tx_data), .C(_91_), .D(_99_), .Y(_7_) );
	INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_1_), .Y(_125_) );
	NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_125_), .Y(_126_) );
	NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_126_), .Y(_127_) );
	NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_98_), .C(_125_), .Y(_128_) );
	OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_0_), .B(tx_cnt_1_), .C(tx_cnt_2_), .Y(_129_) );
	NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_129_), .C(_128_), .Y(_130_) );
	OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_0_), .B(tx_cnt_1_), .C(_98_), .Y(_131_) );
	NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_2_), .B(_86_), .C(_125_), .Y(_132_) );
	OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_3_), .B(tx_cnt_2_), .C(tx_reg_7_), .Y(_133_) );
	NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_133_), .C(_132_), .Y(_134_) );
	NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_134_), .C(_130_), .Y(_135_) );
	NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_129_), .C(_128_), .Y(_136_) );
	NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_2_), .B(_118_), .Y(_137_) );
	NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_137_), .C(_136_), .Y(_138_) );
	NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_138_), .C(_135_), .Y(_139_) );
	NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_129_), .C(_128_), .Y(_140_) );
	OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_3_), .B(tx_cnt_2_), .C(tx_reg_6_), .Y(_141_) );
	NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_141_), .C(_132_), .Y(_142_) );
	NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_142_), .C(_140_), .Y(_143_) );
	NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_129_), .C(_128_), .Y(_144_) );
	NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_2_), .B(_116_), .Y(_145_) );
	NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_145_), .C(_144_), .Y(_146_) );
	NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_0_), .B(_146_), .C(_143_), .Y(_147_) );
	NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_3_), .B(_128_), .Y(_148_) );
	OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(tx_cnt_2_), .B(_126_), .C(tx_cnt_3_), .Y(_149_) );
	NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_149_), .Y(_150_) );
	NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_150_), .Y(_151_) );
	NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_139_), .C(_147_), .Y(_152_) );
	NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_99_), .Y(_153_) );
	AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_170_), .C(_153_), .Y(_154_) );
	NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_152_), .Y(_8_) );
	NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_12_), .Y(_155_) );
	NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_155_), .Y(_156_) );
	MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_163_), .S(_156_), .Y(_4__7_) );
	MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_163_), .S(_53_), .Y(_4__6_) );
	NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_34_), .C(_21_), .Y(_157_) );
	NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(rx_reg_5_), .B(_157_), .Y(_158_) );
	OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_157_), .C(_158_), .Y(_4__5_) );
	OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(rx_busy), .B(_163_), .C(_50_), .Y(_159_) );
	AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(rx_busy), .Y(_160_) );
	OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_44_), .C(_160_), .Y(_161_) );
	AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_159_), .C(_16_), .Y(_0_) );
	INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(_162_) );
	BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_167__0_), .Y(rx_data[0]) );
	BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_167__1_), .Y(rx_data[1]) );
	BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_167__2_), .Y(rx_data[2]) );
	BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_167__3_), .Y(rx_data[3]) );
	BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_167__4_), .Y(rx_data[4]) );
	BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_167__5_), .Y(rx_data[5]) );
	BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_167__6_), .Y(rx_data[6]) );
	BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_167__7_), .Y(rx_data[7]) );
	BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_168_), .Y(rx_empty) );
	BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_169_), .Y(tx_empty) );
	BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_170_), .Y(tx_out) );
	DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_8_), .Q(_170_), .R(vdd), .S(_162__bF_buf5) );
	DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_7_), .Q(_169_), .R(vdd), .S(_162__bF_buf4) );
	DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_9__0_), .Q(tx_reg_0_), .R(_162__bF_buf3), .S(vdd) );
	DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_9__1_), .Q(tx_reg_1_), .R(_162__bF_buf2), .S(vdd) );
	DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_9__2_), .Q(tx_reg_2_), .R(_162__bF_buf1), .S(vdd) );
	DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_9__3_), .Q(tx_reg_3_), .R(_162__bF_buf0), .S(vdd) );
	DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_9__4_), .Q(tx_reg_4_), .R(_162__bF_buf5), .S(vdd) );
	DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_9__5_), .Q(tx_reg_5_), .R(_162__bF_buf4), .S(vdd) );
	DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_9__6_), .Q(tx_reg_6_), .R(_162__bF_buf3), .S(vdd) );
	DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_9__7_), .Q(tx_reg_7_), .R(_162__bF_buf2), .S(vdd) );
	DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_6__0_), .Q(tx_cnt_0_), .R(_162__bF_buf1), .S(vdd) );
	DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_6__1_), .Q(tx_cnt_1_), .R(_162__bF_buf0), .S(vdd) );
	DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_6__2_), .Q(tx_cnt_2_), .R(_162__bF_buf5), .S(vdd) );
	DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(txclk), .D(_6__3_), .Q(tx_cnt_3_), .R(_162__bF_buf4), .S(vdd) );
	DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf4), .D(_2__0_), .Q(_167__0_), .R(_162__bF_buf3), .S(vdd) );
	DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf3), .D(_2__1_), .Q(_167__1_), .R(_162__bF_buf2), .S(vdd) );
	DFFSR DFFSR_17 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf2), .D(_2__2_), .Q(_167__2_), .R(_162__bF_buf1), .S(vdd) );
	DFFSR DFFSR_18 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf1), .D(_2__3_), .Q(_167__3_), .R(_162__bF_buf0), .S(vdd) );
	DFFSR DFFSR_19 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf0), .D(_2__4_), .Q(_167__4_), .R(_162__bF_buf5), .S(vdd) );
	DFFSR DFFSR_20 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf4), .D(_2__5_), .Q(_167__5_), .R(_162__bF_buf4), .S(vdd) );
	DFFSR DFFSR_21 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf3), .D(_2__6_), .Q(_167__6_), .R(_162__bF_buf3), .S(vdd) );
	DFFSR DFFSR_22 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf2), .D(_2__7_), .Q(_167__7_), .R(_162__bF_buf2), .S(vdd) );
	DFFSR DFFSR_23 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf1), .D(_3_), .Q(_168_), .R(vdd), .S(_162__bF_buf1) );
	DFFSR DFFSR_24 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf0), .D(_4__0_), .Q(rx_reg_0_), .R(_162__bF_buf0), .S(vdd) );
	DFFSR DFFSR_25 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf4), .D(_4__1_), .Q(rx_reg_1_), .R(_162__bF_buf5), .S(vdd) );
	DFFSR DFFSR_26 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf3), .D(_4__2_), .Q(rx_reg_2_), .R(_162__bF_buf4), .S(vdd) );
	DFFSR DFFSR_27 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf2), .D(_4__3_), .Q(rx_reg_3_), .R(_162__bF_buf3), .S(vdd) );
	DFFSR DFFSR_28 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf1), .D(_4__4_), .Q(rx_reg_4_), .R(_162__bF_buf2), .S(vdd) );
	DFFSR DFFSR_29 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf0), .D(_4__5_), .Q(rx_reg_5_), .R(_162__bF_buf1), .S(vdd) );
	DFFSR DFFSR_30 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf4), .D(_4__6_), .Q(rx_reg_6_), .R(_162__bF_buf0), .S(vdd) );
	DFFSR DFFSR_31 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf3), .D(_4__7_), .Q(rx_reg_7_), .R(_162__bF_buf5), .S(vdd) );
	DFFSR DFFSR_32 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf2), .D(_5__0_), .Q(rx_sample_cnt_0_), .R(_162__bF_buf4), .S(vdd) );
	DFFSR DFFSR_33 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf1), .D(_5__1_), .Q(rx_sample_cnt_1_), .R(_162__bF_buf3), .S(vdd) );
	DFFSR DFFSR_34 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf0), .D(_5__2_), .Q(rx_sample_cnt_2_), .R(_162__bF_buf2), .S(vdd) );
	DFFSR DFFSR_35 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf4), .D(_5__3_), .Q(rx_sample_cnt_3_), .R(_162__bF_buf1), .S(vdd) );
	DFFSR DFFSR_36 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf3), .D(_1__0_), .Q(rx_cnt_0_), .R(_162__bF_buf0), .S(vdd) );
	DFFSR DFFSR_37 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf2), .D(_1__1_), .Q(rx_cnt_1_), .R(_162__bF_buf5), .S(vdd) );
	DFFSR DFFSR_38 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf1), .D(_1__2_), .Q(rx_cnt_2_), .R(_162__bF_buf4), .S(vdd) );
	DFFSR DFFSR_39 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf0), .D(_1__3_), .Q(rx_cnt_3_), .R(_162__bF_buf3), .S(vdd) );
	DFFSR DFFSR_40 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf4), .D(rx_in), .Q(rx_d1), .R(vdd), .S(_162__bF_buf2) );
	DFFSR DFFSR_41 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf3), .D(rx_d1), .Q(rx_d2), .R(vdd), .S(_162__bF_buf1) );
	DFFSR DFFSR_42 ( .gnd(gnd), .vdd(vdd), .CLK(rxclk_bF_buf2), .D(_0_), .Q(rx_busy), .R(_162__bF_buf0), .S(vdd) );
endmodule
