module counter_b4 (b4_enable, b4_clk, b4_reset, b4_mode, b4_D, b4_load, b4_rco, b4_Q);

input b4_enable;
input b4_clk;
input b4_reset;
output b4_load;
output b4_rco;
input [1:0] b4_mode;
input [3:0] b4_D;
output [3:0] b4_Q;

wire vdd = 1'b1;
wire gnd = 1'b0;

	AOI21X1 AOI21X1_1 ( .A(_38_), .B(_25_), .C(_41_), .Y(_42_) );
	INVX1 INVX1_1 ( .A(b4_D[3]), .Y(_43_) );
	OAI21X1 OAI21X1_1 ( .A(_43_), .B(_8_), .C(_5_), .Y(_44_) );
	AOI21X1 AOI21X1_2 ( .A(_40_), .B(_42_), .C(_44_), .Y(_45_) );
	NAND3X1 NAND3X1_1 ( .A(_23_), .B(_38_), .C(_15_), .Y(_46_) );
	OR2X2 OR2X2_1 ( .A(_56__0_), .B(_56__1_), .Y(_47_) );
	OAI21X1 OAI21X1_2 ( .A(_56__2_), .B(_47_), .C(_56__3_), .Y(_48_) );
	NAND2X1 NAND2X1_1 ( .A(_46_), .B(_48_), .Y(_49_) );
	XNOR2X1 XNOR2X1_1 ( .A(_27_), .B(_38_), .Y(_50_) );
	AOI22X1 AOI22X1_1 ( .A(_24_), .B(_50_), .C(_19_), .D(_49_), .Y(_51_) );
	AOI22X1 AOI22X1_2 ( .A(_38_), .B(_6_), .C(_45_), .D(_51_), .Y(_3__3_) );
	NOR2X1 NOR2X1_1 ( .A(_16_), .B(_6_), .Y(_0__0_) );
	NOR2X1 NOR2X1_2 ( .A(_13_), .B(_6_), .Y(_0__1_) );
	NOR2X1 NOR2X1_3 ( .A(_23_), .B(_6_), .Y(_0__2_) );
	NOR2X1 NOR2X1_4 ( .A(_38_), .B(_6_), .Y(_0__3_) );
	INVX1 INVX1_2 ( .A(_46_), .Y(_52_) );
	NAND2X1 NAND2X1_2 ( .A(_19_), .B(_52_), .Y(_53_) );
	AND2X2 AND2X2_1 ( .A(_27_), .B(_38_), .Y(_54_) );
	AOI22X1 AOI22X1_3 ( .A(_32_), .B(_39_), .C(_24_), .D(_54_), .Y(_55_) );
	AOI21X1 AOI21X1_3 ( .A(_53_), .B(_55_), .C(_6_), .Y(_2_) );
	NOR2X1 NOR2X1_5 ( .A(_8_), .B(_6_), .Y(_1_) );
	BUFX2 BUFX2_1 ( .A(_56__0_), .Y(b4_Q[0]) );
	BUFX2 BUFX2_2 ( .A(_56__1_), .Y(b4_Q[1]) );
	BUFX2 BUFX2_3 ( .A(_56__2_), .Y(b4_Q[2]) );
	BUFX2 BUFX2_4 ( .A(_56__3_), .Y(b4_Q[3]) );
	BUFX2 BUFX2_5 ( .A(_57_), .Y(b4_load) );
	BUFX2 BUFX2_6 ( .A(_58_), .Y(b4_rco) );
	DFFPOSX1 DFFPOSX1_1 ( .CLK(b4_clk), .D(_1_), .Q(_57_) );
	DFFPOSX1 DFFPOSX1_2 ( .CLK(b4_clk), .D(_2_), .Q(_58_) );
	DFFPOSX1 DFFPOSX1_3 ( .CLK(b4_clk), .D(_0__0_), .Q(_56__0_) );
	DFFPOSX1 DFFPOSX1_4 ( .CLK(b4_clk), .D(_0__1_), .Q(_56__1_) );
	DFFPOSX1 DFFPOSX1_5 ( .CLK(b4_clk), .D(_0__2_), .Q(_56__2_) );
	DFFPOSX1 DFFPOSX1_6 ( .CLK(b4_clk), .D(_0__3_), .Q(_56__3_) );
	DFFPOSX1 DFFPOSX1_7 ( .CLK(b4_clk), .D(_3__0_), .Q(_56__0_) );
	DFFPOSX1 DFFPOSX1_8 ( .CLK(b4_clk), .D(_3__1_), .Q(_56__1_) );
	DFFPOSX1 DFFPOSX1_9 ( .CLK(b4_clk), .D(_3__2_), .Q(_56__2_) );
	DFFPOSX1 DFFPOSX1_10 ( .CLK(b4_clk), .D(_3__3_), .Q(_56__3_) );
	INVX1 INVX1_3 ( .A(b4_enable), .Y(_4_) );
	NOR2X1 NOR2X1_6 ( .A(b4_reset), .B(_4_), .Y(_5_) );
	INVX4 INVX4_1 ( .A(_5_), .Y(_6_) );
	OAI21X1 OAI21X1_3 ( .A(b4_reset), .B(_4_), .C(_56__0_), .Y(_7_) );
	NAND2X1 NAND2X1_3 ( .A(b4_mode[0]), .B(b4_mode[1]), .Y(_8_) );
	INVX1 INVX1_4 ( .A(b4_mode[0]), .Y(_9_) );
	INVX1 INVX1_5 ( .A(b4_mode[1]), .Y(_10_) );
	OAI21X1 OAI21X1_4 ( .A(_9_), .B(_10_), .C(_56__0_), .Y(_11_) );
	OAI21X1 OAI21X1_5 ( .A(b4_D[0]), .B(_8_), .C(_11_), .Y(_12_) );
	OAI21X1 OAI21X1_6 ( .A(_6_), .B(_12_), .C(_7_), .Y(_3__0_) );
	INVX1 INVX1_6 ( .A(_56__1_), .Y(_13_) );
	INVX1 INVX1_7 ( .A(_8_), .Y(_14_) );
	NOR2X1 NOR2X1_7 ( .A(_56__0_), .B(_56__1_), .Y(_15_) );
	INVX1 INVX1_8 ( .A(_56__0_), .Y(_16_) );
	NOR2X1 NOR2X1_8 ( .A(_16_), .B(_13_), .Y(_17_) );
	OR2X2 OR2X2_2 ( .A(_17_), .B(_15_), .Y(_18_) );
	NOR2X1 NOR2X1_9 ( .A(b4_mode[1]), .B(_9_), .Y(_19_) );
	AOI22X1 AOI22X1_4 ( .A(b4_D[1]), .B(_14_), .C(_19_), .D(_18_), .Y(_20_) );
	NOR2X1 NOR2X1_10 ( .A(_15_), .B(_17_), .Y(_21_) );
	AOI21X1 AOI21X1_4 ( .A(_21_), .B(_9_), .C(_6_), .Y(_22_) );
	AOI22X1 AOI22X1_5 ( .A(_13_), .B(_6_), .C(_22_), .D(_20_), .Y(_3__1_) );
	INVX2 INVX2_1 ( .A(_56__2_), .Y(_23_) );
	NOR2X1 NOR2X1_11 ( .A(b4_mode[0]), .B(_10_), .Y(_24_) );
	NAND3X1 NAND3X1_2 ( .A(_56__0_), .B(_56__1_), .C(_56__2_), .Y(_25_) );
	INVX1 INVX1_9 ( .A(_25_), .Y(_26_) );
	AOI21X1 AOI21X1_5 ( .A(_56__0_), .B(_56__1_), .C(_56__2_), .Y(_27_) );
	OR2X2 OR2X2_3 ( .A(_26_), .B(_27_), .Y(_28_) );
	INVX1 INVX1_10 ( .A(b4_D[2]), .Y(_29_) );
	OAI21X1 OAI21X1_7 ( .A(_29_), .B(_8_), .C(_5_), .Y(_30_) );
	AOI21X1 AOI21X1_6 ( .A(_28_), .B(_24_), .C(_30_), .Y(_31_) );
	NOR2X1 NOR2X1_12 ( .A(b4_mode[0]), .B(b4_mode[1]), .Y(_32_) );
	NOR2X1 NOR2X1_13 ( .A(_27_), .B(_26_), .Y(_33_) );
	NAND2X1 NAND2X1_4 ( .A(_23_), .B(_15_), .Y(_34_) );
	OAI21X1 OAI21X1_8 ( .A(_56__0_), .B(_56__1_), .C(_56__2_), .Y(_35_) );
	NAND2X1 NAND2X1_5 ( .A(_35_), .B(_34_), .Y(_36_) );
	AOI22X1 AOI22X1_6 ( .A(_36_), .B(_19_), .C(_32_), .D(_33_), .Y(_37_) );
	AOI22X1 AOI22X1_7 ( .A(_23_), .B(_6_), .C(_37_), .D(_31_), .Y(_3__2_) );
	INVX4 INVX4_2 ( .A(_56__3_), .Y(_38_) );
	NOR2X1 NOR2X1_14 ( .A(_38_), .B(_25_), .Y(_39_) );
	INVX1 INVX1_11 ( .A(_39_), .Y(_40_) );
	INVX1 INVX1_12 ( .A(_32_), .Y(_41_) );
endmodule
