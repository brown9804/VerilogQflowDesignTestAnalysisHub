*** SPICE deck for cell NAND3{lay} from library Design_NOR3_NAND3_AOI22
*** Created on Sun Dec 06, 2020 16:40:26
*** Last revised on Sun Dec 06, 2020 17:34:11
*** Written on Sun Dec 06, 2020 18:45:06 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

*** TOP LEVEL CELL: NAND3{lay}
Mnmos@0 net@21 A gnd gnd NMOS L=0.2U W=1.8U AS=2.58P AD=0.54P PS=11.8U PD=2.4U
Mnmos@1 net@26 B net@21 gnd NMOS L=0.2U W=1.8U AS=0.54P AD=0.45P PS=2.4U PD=2.3U
Mnmos@2 A_nand_B_nand_C C net@26 gnd NMOS L=0.2U W=1.8U AS=0.45P AD=0.758P PS=2.3U PD=3.35U
Mpmos@0 vdd A A_nand_B_nand_C vdd PMOS L=0.2U W=1.5U AS=0.758P AD=1.233P PS=3.35U PD=5.533U
Mpmos@1 A_nand_B_nand_C B vdd vdd PMOS L=0.2U W=1.5U AS=1.233P AD=0.758P PS=5.533U PD=3.35U
Mpmos@2 vdd C A_nand_B_nand_C vdd PMOS L=0.2U W=1.5U AS=0.758P AD=1.233P PS=3.35U PD=5.533U
.END
