module counter_b4 ( gnd, vdd, b4_enable, b4_clk, b4_reset, b4_mode, b4_D, b4_load, b4_rco, b4_Q);

input gnd, vdd;
input b4_enable;
input b4_clk;
input b4_reset;
output b4_load;
output b4_rco;
input [1:0] b4_mode;
input [3:0] b4_D;
output [3:0] b4_Q;

	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_5_), .Y(_0__1_) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_5_), .Y(_0__2_) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_5_), .Y(_0__3_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_5_), .Y(_1_) );
	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_48__0_), .Y(b4_Q[0]) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_48__1_), .Y(b4_Q[1]) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_48__2_), .Y(b4_Q[2]) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_48__3_), .Y(b4_Q[3]) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(b4_load) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(b4_rco) );
	DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(b4_clk), .D(_1_), .Q(_49_) );
	DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(b4_clk), .D(_0__0_), .Q(_48__0_) );
	DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(b4_clk), .D(_0__1_), .Q(_48__1_) );
	DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(b4_clk), .D(_0__2_), .Q(_48__2_) );
	DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(b4_clk), .D(_0__3_), .Q(_48__3_) );
	DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(b4_clk), .D(_2__0_), .Q(_48__0_) );
	DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(b4_clk), .D(_2__1_), .Q(_48__1_) );
	DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(b4_clk), .D(_2__2_), .Q(_48__2_) );
	DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(b4_clk), .D(_2__3_), .Q(_48__3_) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(b4_enable), .Y(_3_) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(b4_reset), .B(_3_), .Y(_4_) );
	INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_5_) );
	OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(b4_reset), .B(_3_), .C(_48__0_), .Y(_6_) );
	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(b4_mode[0]), .B(b4_mode[1]), .Y(_7_) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(b4_mode[0]), .Y(_8_) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(b4_mode[1]), .Y(_9_) );
	OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_9_), .C(_48__0_), .Y(_10_) );
	OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(b4_D[0]), .B(_7_), .C(_10_), .Y(_11_) );
	OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_11_), .C(_6_), .Y(_2__0_) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_48__1_), .Y(_12_) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_48__0_), .Y(_13_) );
	NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_12_), .Y(_14_) );
	NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_48__0_), .B(_48__1_), .Y(_15_) );
	OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_15_), .Y(_16_) );
	OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(b4_mode[0]), .Y(_17_) );
	NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(b4_mode[1]), .B(_8_), .Y(_18_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(b4_D[1]), .Y(_19_) );
	OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_7_), .C(_4_), .Y(_20_) );
	AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_18_), .C(_20_), .Y(_21_) );
	AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_5_), .C(_21_), .D(_17_), .Y(_2__1_) );
	INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(_48__2_), .Y(_22_) );
	NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(b4_mode[0]), .B(b4_mode[1]), .Y(_23_) );
	NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_48__0_), .B(_48__1_), .C(_48__2_), .Y(_24_) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_24_), .Y(_25_) );
	AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_48__0_), .B(_48__1_), .C(_48__2_), .Y(_26_) );
	NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_25_), .Y(_27_) );
	INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(b4_D[2]), .Y(_28_) );
	OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_7_), .C(_4_), .Y(_29_) );
	AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_23_), .C(_29_), .Y(_30_) );
	XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_22_), .Y(_31_) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(b4_mode[1]), .B(_8_), .Y(_32_) );
	INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_26_), .Y(_33_) );
	AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_24_), .C(_32_), .Y(_34_) );
	AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_18_), .C(_34_), .Y(_35_) );
	AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_5_), .C(_30_), .D(_35_), .Y(_2__2_) );
	INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(_48__3_), .Y(_36_) );
	INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_23_), .Y(_37_) );
	OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_26_), .C(_37_), .D(_25_), .Y(_38_) );
	INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(b4_D[3]), .Y(_39_) );
	OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_7_), .C(_4_), .Y(_40_) );
	AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_48__3_), .C(_40_), .Y(_41_) );
	OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_48__0_), .B(_48__1_), .Y(_42_) );
	OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_48__2_), .B(_42_), .C(_48__3_), .Y(_43_) );
	NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_36_), .C(_15_), .Y(_44_) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_43_), .Y(_45_) );
	OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_24_), .C(_32_), .D(_33_), .Y(_46_) );
	AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_46_), .C(_18_), .D(_45_), .Y(_47_) );
	AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_5_), .C(_41_), .D(_47_), .Y(_2__3_) );
	NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_5_), .Y(_0__0_) );
endmodule
